module AXI4StreamWidthAdapater_4_to_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [7:0]  auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [7:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg [1:0] _T_3; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire  _T_4; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire  _T_5; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_6; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_7; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_9; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_10; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_12; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_13; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_15; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_16; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [23:0] _T_18; // @[Cat.scala 29:58]
  wire  ov0; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg  _T_20; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_4;
  reg  _T_21; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_5;
  reg  _T_22; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_6;
  reg [1:0] _T_23; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_7;
  wire  _T_25; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_26; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_27; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_29; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_30; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_32; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_33; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_35; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_36; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [3:0] _T_39; // @[Cat.scala 29:58]
  wire  ov1; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_44; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_8;
  wire  _T_46; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_47; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_48; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_8; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_64; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_9;
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_67; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_68; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_12; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_84; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_10;
  wire  _T_86; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_87; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_88; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_16; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_101; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_104; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_105; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_108; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_109; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_112; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_113; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_116; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_4 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  assign _T_5 = _T_3 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_6 = _T_3 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_7 = _T_5 ? 3'h0 : _T_6; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_0 = _T_4 ? _T_7 : {{1'd0}, _T_3}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_9 = _T_3 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_10 = _T_4 & _T_9; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_12 = _T_3 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_13 = _T_4 & _T_12; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_15 = _T_3 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_16 = _T_4 & _T_15; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_18 = {auto_in_bits_data,_T_2,_T_1}; // @[Cat.scala 29:58]
  assign ov0 = _T_5 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_25 = _T_23 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_26 = _T_23 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_27 = _T_25 ? 3'h0 : _T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_4 = _T_4 ? _T_27 : {{1'd0}, _T_23}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_29 = _T_23 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_30 = _T_4 & _T_29; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_32 = _T_23 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_33 = _T_4 & _T_32; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_35 = _T_23 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_36 = _T_4 & _T_35; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_39 = {auto_in_bits_last,_T_22,_T_21,_T_20}; // @[Cat.scala 29:58]
  assign ov1 = _T_25 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_46 = _T_44 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_47 = _T_44 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_48 = _T_46 ? 3'h0 : _T_47; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_8 = _T_4 ? _T_48 : {{1'd0}, _T_44}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov2 = _T_46 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_66 = _T_64 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_67 = _T_64 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_68 = _T_66 ? 3'h0 : _T_67; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_12 = _T_4 ? _T_68 : {{1'd0}, _T_64}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov3 = _T_66 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_86 = _T_84 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_87 = _T_84 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_88 = _T_86 ? 3'h0 : _T_87; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_16 = _T_4 ? _T_88 : {{1'd0}, _T_84}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov4 = _T_86 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_101 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  assign _T_103 = _T_101 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_104 = ~_T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_105 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  assign _T_107 = _T_105 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_108 = ~_T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_109 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  assign _T_111 = _T_109 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_112 = ~_T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_113 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  assign _T_115 = _T_113 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_116 = ~_T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_5 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {_T_18,_T}; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = _T_39 != 4'h0; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_20 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_23 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_44 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_64 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_84 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_10) begin
      _T <= auto_in_bits_data;
    end
    if (_T_13) begin
      _T_1 <= auto_in_bits_data;
    end
    if (_T_16) begin
      _T_2 <= auto_in_bits_data;
    end
    if (reset) begin
      _T_3 <= 2'h0;
    end else begin
      _T_3 <= _GEN_0[1:0];
    end
    if (_T_30) begin
      _T_20 <= auto_in_bits_last;
    end
    if (_T_33) begin
      _T_21 <= auto_in_bits_last;
    end
    if (_T_36) begin
      _T_22 <= auto_in_bits_last;
    end
    if (reset) begin
      _T_23 <= 2'h0;
    end else begin
      _T_23 <= _GEN_4[1:0];
    end
    if (reset) begin
      _T_44 <= 2'h0;
    end else begin
      _T_44 <= _GEN_8[1:0];
    end
    if (reset) begin
      _T_64 <= 2'h0;
    end else begin
      _T_64 <= _GEN_12[1:0];
    end
    if (reset) begin
      _T_84 <= 2'h0;
    end else begin
      _T_84 <= _GEN_16[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_108) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_108) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_112) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_116) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_116) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_extra
);
  reg  _T_read [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_read__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_read__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_read__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_extra [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire  _T_extra__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_extra__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_read__T_18_addr = value_1;
  assign _T_read__T_18_data = _T_read[_T_read__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_read__T_10_data = io_enq_bits_read;
  assign _T_read__T_10_addr = value;
  assign _T_read__T_10_mask = 1'h1;
  assign _T_read__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_extra__T_18_addr = value_1;
  assign _T_extra__T_18_data = _T_extra[_T_extra__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_extra__T_10_data = io_enq_bits_extra;
  assign _T_extra__T_10_addr = value;
  assign _T_extra__T_10_mask = 1'h1;
  assign _T_extra__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_read = _T_read__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_extra = _T_extra__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_extra[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_read__T_10_en & _T_read__T_10_mask) begin
      _T_read[_T_read__T_10_addr] <= _T_read__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_extra__T_10_en & _T_extra__T_10_mask) begin
      _T_extra[_T_extra__T_10_addr] <= _T_extra__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4Splitter(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_4_ready,
  output        auto_stream_out_4_valid,
  output [31:0] auto_stream_out_4_bits_data,
  output        auto_stream_out_4_bits_last,
  input         auto_stream_out_3_ready,
  output        auto_stream_out_3_valid,
  output [31:0] auto_stream_out_3_bits_data,
  output        auto_stream_out_3_bits_last,
  input         auto_stream_out_2_ready,
  output        auto_stream_out_2_valid,
  output [31:0] auto_stream_out_2_bits_data,
  output        auto_stream_out_2_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_7; // @[RegisterRouter.scala 40:39]
  wire  _T_8; // @[RegisterRouter.scala 40:26]
  wire  _T_9; // @[RegisterRouter.scala 42:29]
  wire  _T_52_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_16; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_56; // @[RegisterRouter.scala 59:16]
  wire  _T_58; // @[RegisterRouter.scala 59:16]
  wire  _T_10; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_19; // @[OneHot.scala 65:12]
  wire [1:0] _T_21; // @[Misc.scala 200:81]
  wire  _T_22; // @[Misc.scala 204:21]
  wire  _T_25; // @[Misc.scala 209:20]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_30; // @[Misc.scala 213:38]
  wire  _T_31; // @[Misc.scala 213:29]
  wire  _T_34; // @[Misc.scala 209:20]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 212:27]
  wire  _T_45; // @[Misc.scala 213:38]
  wire  _T_46; // @[Misc.scala 213:29]
  wire [3:0] _T_49; // @[Cat.scala 29:58]
  wire [3:0] _T_51; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_70; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76; // @[Bitwise.scala 72:12]
  wire [31:0] _T_79; // @[Cat.scala 29:58]
  wire  _T_98; // @[RegisterRouter.scala 59:16]
  wire  _T_151; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_145; // @[OneHot.scala 58:35]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_175; // @[RegisterRouter.scala 59:16]
  wire  _T_176; // @[RegisterRouter.scala 59:16]
  wire  _T_105; // @[RegisterRouter.scala 59:16]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_171; // @[RegisterRouter.scala 59:16]
  wire  _T_128; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_226_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_226_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_229; // @[RegisterRouter.scala 65:29]
  wire  _T_232; // @[Splitter.scala 45:34]
  wire  _T_233; // @[Splitter.scala 45:34]
  wire  _T_234; // @[Splitter.scala 45:34]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  _T_235; // @[Splitter.scala 46:34]
  wire  _T_236; // @[Splitter.scala 46:34]
  wire  _T_237; // @[Splitter.scala 46:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_238; // @[Splitter.scala 49:19]
  wire  _T_239; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_242; // @[Splitter.scala 62:34]
  wire  _T_246; // @[Splitter.scala 62:34]
  wire  _T_250; // @[Splitter.scala 62:34]
  wire  _T_254; // @[Splitter.scala 62:34]
  wire  _T_258; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_7 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_8 = auto_mem_in_ar_valid | _T_7; // @[RegisterRouter.scala 40:26]
  assign _T_9 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_52_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_16 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_56 = _T_16[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_58 = _T_56 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_10 = _T_52_ready & _T_9; // @[RegisterRouter.scala 42:26]
  assign _T_19 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_21 = _T_19 | 2'h1; // @[Misc.scala 200:81]
  assign _T_22 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_25 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_27 = _T_21[1] & _T_25; // @[Misc.scala 213:38]
  assign _T_28 = _T_22 | _T_27; // @[Misc.scala 213:29]
  assign _T_30 = _T_21[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_31 = _T_22 | _T_30; // @[Misc.scala 213:29]
  assign _T_34 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_35 = _T_25 & _T_34; // @[Misc.scala 212:27]
  assign _T_36 = _T_21[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = _T_25 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_39 = _T_21[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & _T_34; // @[Misc.scala 212:27]
  assign _T_42 = _T_21[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_31 | _T_42; // @[Misc.scala 213:29]
  assign _T_44 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_45 = _T_21[0] & _T_44; // @[Misc.scala 213:38]
  assign _T_46 = _T_31 | _T_45; // @[Misc.scala 213:29]
  assign _T_49 = {_T_46,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  assign _T_51 = auto_mem_in_ar_valid ? _T_49 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_70 = _T_51[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_72 = _T_51[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_74 = _T_51[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = _T_51[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_79 = {_T_76,_T_74,_T_72,_T_70}; // @[Cat.scala 29:58]
  assign _T_98 = _T_79 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_151 = _T_8 & _T_52_ready; // @[RegisterRouter.scala 59:16]
  assign _T_145 = 2'h1 << _T_16[2]; // @[OneHot.scala 58:35]
  assign _T_168 = _T_151 & _T_9; // @[RegisterRouter.scala 59:16]
  assign _T_175 = _T_168 & _T_145[1]; // @[RegisterRouter.scala 59:16]
  assign _T_176 = _T_175 & _T_58; // @[RegisterRouter.scala 59:16]
  assign _T_105 = _T_176 & _T_98; // @[RegisterRouter.scala 59:16]
  assign _T_170 = _T_168 & _T_145[0]; // @[RegisterRouter.scala 59:16]
  assign _T_171 = _T_170 & _T_58; // @[RegisterRouter.scala 59:16]
  assign _T_128 = _T_171 & _T_98; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_16[2] ? _T_58 : _T_58; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_16[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_226_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_226_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_229 = ~_T_226_bits_read; // @[RegisterRouter.scala 65:29]
  assign _T_232 = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign _T_233 = _T_232 | auto_stream_out_2_ready; // @[Splitter.scala 45:34]
  assign _T_234 = _T_233 | auto_stream_out_3_ready; // @[Splitter.scala 45:34]
  assign readyOR = _T_234 | auto_stream_out_4_ready; // @[Splitter.scala 45:34]
  assign _T_235 = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_236 = _T_235 & auto_stream_out_2_ready; // @[Splitter.scala 46:34]
  assign _T_237 = _T_236 & auto_stream_out_3_ready; // @[Splitter.scala 46:34]
  assign readyAND = _T_237 & auto_stream_out_4_ready; // @[Splitter.scala 46:34]
  assign _T_238 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_239 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_239 & readyOR; // @[Splitter.scala 52:33]
  assign _T_242 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_246 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign _T_250 = ~maskReg[2]; // @[Splitter.scala 62:34]
  assign _T_254 = ~maskReg[3]; // @[Splitter.scala 62:34]
  assign _T_258 = ~maskReg[4]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_10 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_10 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_226_valid & _T_229; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_226_valid & _T_226_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_238 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_4_valid = auto_stream_in_valid & _T_258; // @[LazyModule.scala 173:49]
  assign auto_stream_out_4_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_4_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_valid = auto_stream_in_valid & _T_254; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_valid = auto_stream_in_valid & _T_250; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_246; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_242; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_7; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_226_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_128) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_105) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module Queue_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits_data,
  input        io_enq_bits_last,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits_data,
  output       io_deq_bits_last
);
  reg [7:0] _T_data [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T_data__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 209:24]
  wire [7:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[Decoupled.scala 240:27]
  wire  _GEN_22; // @[Decoupled.scala 237:18]
  wire  _GEN_21; // @[Decoupled.scala 237:18]
  wire  _T_11; // @[Decoupled.scala 227:16]
  wire  _T_12; // @[Decoupled.scala 231:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 237:18]
  assign _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 227:16]
  assign _T_12 = ~_T_3; // @[Decoupled.scala 231:19]
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer(
  input        clock,
  input        reset,
  input        auto_out_out_ready,
  output       auto_out_out_valid,
  output [7:0] auto_out_out_bits_data,
  output       auto_out_out_bits_last,
  output       auto_in_in_ready,
  input        auto_in_in_valid,
  input  [7:0] auto_in_in_bits_data,
  input        auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [7:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [7:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_1 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module PEControlLogic(
  input   io_currCompOut,
  input   io_leftCompOut,
  input   io_rightCompOut,
  input   io_currDiscard,
  input   io_rightPropDiscard,
  output  io_propDiscard,
  output  io_load,
  output  io_leftRightShift,
  output  io_rstPEregs
);
  wire  _T; // @[ControlLogic.scala 24:27]
  wire  load; // @[ControlLogic.scala 24:50]
  wire  _T_4; // @[ControlLogic.scala 30:45]
  wire  _T_5; // @[ControlLogic.scala 30:43]
  wire  _T_6; // @[ControlLogic.scala 30:65]
  wire  _T_7; // @[ControlLogic.scala 30:82]
  wire  _T_9; // @[ControlLogic.scala 30:62]
  assign _T = io_currCompOut ^ io_rightPropDiscard; // @[ControlLogic.scala 24:27]
  assign load = _T | io_currDiscard; // @[ControlLogic.scala 24:50]
  assign _T_4 = ~io_currCompOut; // @[ControlLogic.scala 30:45]
  assign _T_5 = io_leftCompOut & _T_4; // @[ControlLogic.scala 30:43]
  assign _T_6 = ~io_rightCompOut; // @[ControlLogic.scala 30:65]
  assign _T_7 = _T_6 & io_currCompOut; // @[ControlLogic.scala 30:82]
  assign _T_9 = _T_5 + _T_7; // @[ControlLogic.scala 30:62]
  assign io_propDiscard = io_currDiscard | io_rightPropDiscard; // @[ControlLogic.scala 28:18]
  assign io_load = _T | io_currDiscard; // @[ControlLogic.scala 26:11]
  assign io_leftRightShift = io_currCompOut & load; // @[ControlLogic.scala 27:21]
  assign io_rstPEregs = load & _T_9; // @[ControlLogic.scala 30:16]
endmodule
module PE(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_rightOutData,
  output        io_currDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign rightOrLeftCNT = io_lastCell ? 5'h0 : io_rightNBR_lifeCNT; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_rightOutData = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = 1'h1; // @[PE.scala 56:30]
  assign ctrlLogic_io_rightCompOut = _T_3 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_3 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= 16'sh0;
      end else begin
        saveCellData <= io_rightNBR_data;
      end
    end
    if (reset) begin
      cntLife <= 5'h0;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_1(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h1; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h1;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_2(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h2; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h2;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_3(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h3; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h3;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_4(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h4; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h4;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_5(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h5; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h5;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_6(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h6; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h6;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_7(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h7; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h7;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_8(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h8; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h8;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_9(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h9; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h9;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_10(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'ha; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'ha;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_11(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'hb; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'hb;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_12(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'hc; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'hc;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_13(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'hd; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'hd;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_14(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'he; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'he;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_15(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'hf; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'hf;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_16(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h10; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h10;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_17(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h11; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h11;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_18(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h12; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h12;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_19(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h13; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h13;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_20(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h14; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h14;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_21(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h15; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h15;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_22(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input  [4:0]  io_rightNBR_lifeCNT,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? io_rightNBR_lifeCNT : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h16; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h16;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module PE_23(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input  [4:0]  io_leftNBR_lifeCNT,
  input         io_leftNBR_compRes,
  output [15:0] io_currCell_data,
  output [4:0]  io_currCell_lifeCNT,
  output        io_currCell_compRes,
  input  [5:0]  io_lisSize,
  input         io_lastCell,
  input         io_active,
  input  [15:0] io_inData,
  output [15:0] io_leftOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  load; // @[PE.scala 89:29]
  wire [4:0] _T_8; // @[PE.scala 99:26]
  wire [4:0] _GEN_3; // @[PE.scala 97:61]
  wire [4:0] rightOrLeftCNT; // @[PE.scala 93:65]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  reg [4:0] cntLife; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_1;
  wire [5:0] _T_13; // @[LISutil.scala 38:39]
  wire [5:0] _GEN_13; // @[LISutil.scala 38:23]
  wire  discard; // @[LISutil.scala 38:23]
  wire [4:0] _T_15; // @[LISutil.scala 46:44]
  wire [4:0] _T_17; // @[LISutil.scala 41:22]
  wire  _T_18; // @[LISutil.scala 55:17]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_8 = ctrlLogic_io_leftRightShift ? 5'h0 : io_leftNBR_lifeCNT; // @[PE.scala 99:26]
  assign _GEN_3 = io_active ? _T_8 : 5'h17; // @[PE.scala 97:61]
  assign rightOrLeftCNT = io_lastCell ? io_leftNBR_lifeCNT : _GEN_3; // @[PE.scala 93:65]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_13 = io_lisSize - 6'h1; // @[LISutil.scala 38:39]
  assign _GEN_13 = {{1'd0}, cntLife}; // @[LISutil.scala 38:23]
  assign discard = _GEN_13 == _T_13; // @[LISutil.scala 38:23]
  assign _T_15 = rightOrLeftCNT + 5'h1; // @[LISutil.scala 46:44]
  assign _T_17 = cntLife + 5'h1; // @[LISutil.scala 41:22]
  assign _T_18 = ctrlLogic_io_rstPEregs & io_enableSort; // @[LISutil.scala 55:17]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_lifeCNT = cntLife; // @[PE.scala 164:25]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 163:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = 1'h0; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = _GEN_13 == _T_13; // @[PE.scala 162:30]
  assign ctrlLogic_io_rightPropDiscard = 1'h0; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntLife = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= 16'sh0;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
    if (reset) begin
      cntLife <= 5'h17;
    end else if (_T_18) begin
      cntLife <= 5'h0;
    end else if (load) begin
      cntLife <= _T_15;
    end else if (io_enableSort) begin
      if (discard) begin
        cntLife <= 5'h0;
      end else begin
        cntLife <= _T_17;
      end
    end
  end
endmodule
module LinearSorter(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut,
  output [15:0] io_sortedData_0,
  output [15:0] io_sortedData_1,
  output [15:0] io_sortedData_2,
  output [15:0] io_sortedData_3,
  output [15:0] io_sortedData_4,
  output [15:0] io_sortedData_5,
  output [15:0] io_sortedData_6,
  output [15:0] io_sortedData_7,
  output [15:0] io_sortedData_8,
  output [15:0] io_sortedData_9,
  output [15:0] io_sortedData_10,
  output [15:0] io_sortedData_11,
  output [15:0] io_sortedData_12,
  output [15:0] io_sortedData_13,
  output [15:0] io_sortedData_14,
  output [15:0] io_sortedData_15,
  output [15:0] io_sortedData_16,
  output [15:0] io_sortedData_17,
  output [15:0] io_sortedData_18,
  output [15:0] io_sortedData_19,
  output [15:0] io_sortedData_20,
  output [15:0] io_sortedData_21,
  output [15:0] io_sortedData_22,
  output [15:0] io_sortedData_23,
  output        io_sorterFull,
  output        io_sorterEmpty,
  input  [5:0]  io_lisSize
);
  wire  PEChain_0_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_0_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_0_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_0_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_0_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_lastCell; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_1_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_1_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_1_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_1_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_1_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_2_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_2_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_2_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_2_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_2_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_3_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_3_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_3_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_3_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_3_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_4_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_4_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_4_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_4_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_4_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_5_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_5_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_5_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_5_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_5_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_6_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_6_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_6_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_6_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_6_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_7_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_7_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_7_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_7_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_7_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_8_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_8_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_8_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_8_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_8_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_9_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_9_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_9_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_9_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_9_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_10_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_10_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_10_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_10_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_10_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_11_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_11_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_11_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_11_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_11_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_12_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_12_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_12_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_12_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_12_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_13_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_13_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_13_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_13_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_13_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_14_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_14_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_14_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_14_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_14_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_15_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_15_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_15_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_15_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_15_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_16_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_16_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_16_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_16_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_16_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_17_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_17_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_17_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_17_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_17_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_18_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_18_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_18_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_18_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_18_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_19_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_19_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_19_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_19_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_19_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_20_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_20_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_20_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_20_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_20_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_21_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_21_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_21_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_21_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_21_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_22_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_22_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_22_io_rightNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_22_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_22_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_23_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_23_io_leftNBR_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire [4:0] PEChain_23_io_currCell_lifeCNT; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire [5:0] PEChain_23_io_lisSize; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_active; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_inData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  reg  initialInDone; // @[LinearSorter.scala 67:30]
  reg [31:0] _RAND_0;
  reg [4:0] cntInData; // @[LinearSorter.scala 68:26]
  reg [31:0] _RAND_1;
  reg [1:0] state; // @[LinearSorter.scala 78:22]
  reg [31:0] _RAND_2;
  reg [5:0] lisSizeReg; // @[LinearSorter.scala 81:27]
  reg [31:0] _RAND_3;
  wire [5:0] _T_1; // @[LinearSorter.scala 86:43]
  wire  _T_96; // @[Decoupled.scala 40:37]
  wire [4:0] _T_98; // @[LinearSorter.scala 92:28]
  wire  _T_99; // @[LinearSorter.scala 94:20]
  wire [5:0] _GEN_39; // @[LinearSorter.scala 98:19]
  wire  _T_102; // @[LinearSorter.scala 98:19]
  wire  _T_104; // @[LinearSorter.scala 98:42]
  wire  _T_113; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_7; // @[LinearSorter.scala 117:27]
  wire  _T_115; // @[Conditional.scala 37:30]
  wire  fireLastIn; // @[LinearSorter.scala 111:30]
  wire [1:0] _GEN_8; // @[LinearSorter.scala 120:62]
  wire  _T_117; // @[Conditional.scala 37:30]
  reg [4:0] cntOutData; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_4;
  wire [5:0] _GEN_40; // @[LinearSorter.scala 125:28]
  wire  _T_120; // @[LinearSorter.scala 125:28]
  wire [1:0] _GEN_9; // @[LinearSorter.scala 125:50]
  wire [1:0] _GEN_10; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_11; // @[Conditional.scala 39:67]
  wire [1:0] state_next; // @[Conditional.scala 40:58]
  wire  _T_105; // @[LinearSorter.scala 101:25]
  wire  _GEN_2; // @[LinearSorter.scala 101:36]
  wire  _GEN_3; // @[LinearSorter.scala 98:59]
  wire  _T_106; // @[LinearSorter.scala 106:29]
  wire  _T_107; // @[LinearSorter.scala 106:54]
  wire  enable; // @[LinearSorter.scala 106:45]
  wire  _T_109; // @[LISutil.scala 13:24]
  wire [4:0] _T_111; // @[LISutil.scala 14:22]
  wire  _T_126; // @[LinearSorter.scala 168:63]
  wire  discardSignals_2; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_1; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_0; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_5; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_4; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_3; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [5:0] _T_293; // @[LinearSorter.scala 177:50]
  wire  discardSignals_8; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_7; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_6; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_11; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_10; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_9; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [11:0] _T_299; // @[LinearSorter.scala 177:50]
  wire  discardSignals_14; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_13; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_12; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_17; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_16; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_15; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [5:0] _T_304; // @[LinearSorter.scala 177:50]
  wire  discardSignals_20; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_19; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_18; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_23; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_22; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_21; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [23:0] _T_311; // @[LinearSorter.scala 177:50]
  wire [4:0] _T_336; // @[Mux.scala 47:69]
  wire [4:0] _T_337; // @[Mux.scala 47:69]
  wire [4:0] _T_338; // @[Mux.scala 47:69]
  wire [4:0] _T_339; // @[Mux.scala 47:69]
  wire [4:0] _T_340; // @[Mux.scala 47:69]
  wire [4:0] _T_341; // @[Mux.scala 47:69]
  wire [4:0] _T_342; // @[Mux.scala 47:69]
  wire [4:0] _T_343; // @[Mux.scala 47:69]
  wire [4:0] _T_344; // @[Mux.scala 47:69]
  wire [4:0] _T_345; // @[Mux.scala 47:69]
  wire [4:0] _T_346; // @[Mux.scala 47:69]
  wire [4:0] _T_347; // @[Mux.scala 47:69]
  wire [4:0] _T_348; // @[Mux.scala 47:69]
  wire [4:0] _T_349; // @[Mux.scala 47:69]
  wire [4:0] _T_350; // @[Mux.scala 47:69]
  wire [4:0] _T_351; // @[Mux.scala 47:69]
  wire [4:0] _T_352; // @[Mux.scala 47:69]
  wire [4:0] _T_353; // @[Mux.scala 47:69]
  wire [4:0] _T_354; // @[Mux.scala 47:69]
  wire [4:0] _T_355; // @[Mux.scala 47:69]
  wire [4:0] _T_356; // @[Mux.scala 47:69]
  wire [4:0] _T_357; // @[Mux.scala 47:69]
  wire [4:0] getDiscarded; // @[Mux.scala 47:69]
  wire  _T_359; // @[LinearSorter.scala 199:49]
  wire [15:0] outputData_0; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] outputData_1; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_16; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_2; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_17; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_3; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_18; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_4; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_19; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_5; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_20; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_6; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_21; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_7; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_22; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_8; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_23; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_9; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_24; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_10; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_25; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_11; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_26; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_12; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_27; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_13; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_28; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_14; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_29; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_15; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_30; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_16; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_31; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_17; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_32; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_18; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_33; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_19; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_34; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_20; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_35; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_21; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_36; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_22; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_37; // @[LinearSorter.scala 206:15]
  wire [15:0] outputData_23; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire  _T_365; // @[LinearSorter.scala 208:18]
  wire  _T_367; // @[LinearSorter.scala 208:49]
  wire  _T_369; // @[LinearSorter.scala 209:33]
  PE PEChain_0 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_0_clock),
    .reset(PEChain_0_reset),
    .io_enableSort(PEChain_0_io_enableSort),
    .io_state(PEChain_0_io_state),
    .io_rightNBR_data(PEChain_0_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_0_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_0_io_rightNBR_compRes),
    .io_currCell_data(PEChain_0_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_0_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_0_io_currCell_compRes),
    .io_lisSize(PEChain_0_io_lisSize),
    .io_lastCell(PEChain_0_io_lastCell),
    .io_inData(PEChain_0_io_inData),
    .io_rightPropDiscard(PEChain_0_io_rightPropDiscard),
    .io_rightOutData(PEChain_0_io_rightOutData),
    .io_currDiscard(PEChain_0_io_currDiscard)
  );
  PE_1 PEChain_1 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_1_clock),
    .reset(PEChain_1_reset),
    .io_enableSort(PEChain_1_io_enableSort),
    .io_state(PEChain_1_io_state),
    .io_leftNBR_data(PEChain_1_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_1_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_1_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_1_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_1_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_1_io_rightNBR_compRes),
    .io_currCell_data(PEChain_1_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_1_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_1_io_currCell_compRes),
    .io_lisSize(PEChain_1_io_lisSize),
    .io_lastCell(PEChain_1_io_lastCell),
    .io_active(PEChain_1_io_active),
    .io_inData(PEChain_1_io_inData),
    .io_rightPropDiscard(PEChain_1_io_rightPropDiscard),
    .io_leftOutData(PEChain_1_io_leftOutData),
    .io_rightOutData(PEChain_1_io_rightOutData),
    .io_currDiscard(PEChain_1_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_1_io_toLeftPropDiscard)
  );
  PE_2 PEChain_2 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_2_clock),
    .reset(PEChain_2_reset),
    .io_enableSort(PEChain_2_io_enableSort),
    .io_state(PEChain_2_io_state),
    .io_leftNBR_data(PEChain_2_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_2_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_2_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_2_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_2_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_2_io_rightNBR_compRes),
    .io_currCell_data(PEChain_2_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_2_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_2_io_currCell_compRes),
    .io_lisSize(PEChain_2_io_lisSize),
    .io_lastCell(PEChain_2_io_lastCell),
    .io_active(PEChain_2_io_active),
    .io_inData(PEChain_2_io_inData),
    .io_rightPropDiscard(PEChain_2_io_rightPropDiscard),
    .io_leftOutData(PEChain_2_io_leftOutData),
    .io_rightOutData(PEChain_2_io_rightOutData),
    .io_currDiscard(PEChain_2_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_2_io_toLeftPropDiscard)
  );
  PE_3 PEChain_3 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_3_clock),
    .reset(PEChain_3_reset),
    .io_enableSort(PEChain_3_io_enableSort),
    .io_state(PEChain_3_io_state),
    .io_leftNBR_data(PEChain_3_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_3_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_3_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_3_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_3_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_3_io_rightNBR_compRes),
    .io_currCell_data(PEChain_3_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_3_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_3_io_currCell_compRes),
    .io_lisSize(PEChain_3_io_lisSize),
    .io_lastCell(PEChain_3_io_lastCell),
    .io_active(PEChain_3_io_active),
    .io_inData(PEChain_3_io_inData),
    .io_rightPropDiscard(PEChain_3_io_rightPropDiscard),
    .io_leftOutData(PEChain_3_io_leftOutData),
    .io_rightOutData(PEChain_3_io_rightOutData),
    .io_currDiscard(PEChain_3_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_3_io_toLeftPropDiscard)
  );
  PE_4 PEChain_4 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_4_clock),
    .reset(PEChain_4_reset),
    .io_enableSort(PEChain_4_io_enableSort),
    .io_state(PEChain_4_io_state),
    .io_leftNBR_data(PEChain_4_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_4_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_4_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_4_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_4_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_4_io_rightNBR_compRes),
    .io_currCell_data(PEChain_4_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_4_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_4_io_currCell_compRes),
    .io_lisSize(PEChain_4_io_lisSize),
    .io_lastCell(PEChain_4_io_lastCell),
    .io_active(PEChain_4_io_active),
    .io_inData(PEChain_4_io_inData),
    .io_rightPropDiscard(PEChain_4_io_rightPropDiscard),
    .io_leftOutData(PEChain_4_io_leftOutData),
    .io_rightOutData(PEChain_4_io_rightOutData),
    .io_currDiscard(PEChain_4_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_4_io_toLeftPropDiscard)
  );
  PE_5 PEChain_5 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_5_clock),
    .reset(PEChain_5_reset),
    .io_enableSort(PEChain_5_io_enableSort),
    .io_state(PEChain_5_io_state),
    .io_leftNBR_data(PEChain_5_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_5_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_5_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_5_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_5_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_5_io_rightNBR_compRes),
    .io_currCell_data(PEChain_5_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_5_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_5_io_currCell_compRes),
    .io_lisSize(PEChain_5_io_lisSize),
    .io_lastCell(PEChain_5_io_lastCell),
    .io_active(PEChain_5_io_active),
    .io_inData(PEChain_5_io_inData),
    .io_rightPropDiscard(PEChain_5_io_rightPropDiscard),
    .io_leftOutData(PEChain_5_io_leftOutData),
    .io_rightOutData(PEChain_5_io_rightOutData),
    .io_currDiscard(PEChain_5_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_5_io_toLeftPropDiscard)
  );
  PE_6 PEChain_6 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_6_clock),
    .reset(PEChain_6_reset),
    .io_enableSort(PEChain_6_io_enableSort),
    .io_state(PEChain_6_io_state),
    .io_leftNBR_data(PEChain_6_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_6_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_6_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_6_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_6_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_6_io_rightNBR_compRes),
    .io_currCell_data(PEChain_6_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_6_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_6_io_currCell_compRes),
    .io_lisSize(PEChain_6_io_lisSize),
    .io_lastCell(PEChain_6_io_lastCell),
    .io_active(PEChain_6_io_active),
    .io_inData(PEChain_6_io_inData),
    .io_rightPropDiscard(PEChain_6_io_rightPropDiscard),
    .io_leftOutData(PEChain_6_io_leftOutData),
    .io_rightOutData(PEChain_6_io_rightOutData),
    .io_currDiscard(PEChain_6_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_6_io_toLeftPropDiscard)
  );
  PE_7 PEChain_7 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_7_clock),
    .reset(PEChain_7_reset),
    .io_enableSort(PEChain_7_io_enableSort),
    .io_state(PEChain_7_io_state),
    .io_leftNBR_data(PEChain_7_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_7_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_7_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_7_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_7_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_7_io_rightNBR_compRes),
    .io_currCell_data(PEChain_7_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_7_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_7_io_currCell_compRes),
    .io_lisSize(PEChain_7_io_lisSize),
    .io_lastCell(PEChain_7_io_lastCell),
    .io_active(PEChain_7_io_active),
    .io_inData(PEChain_7_io_inData),
    .io_rightPropDiscard(PEChain_7_io_rightPropDiscard),
    .io_leftOutData(PEChain_7_io_leftOutData),
    .io_rightOutData(PEChain_7_io_rightOutData),
    .io_currDiscard(PEChain_7_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_7_io_toLeftPropDiscard)
  );
  PE_8 PEChain_8 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_8_clock),
    .reset(PEChain_8_reset),
    .io_enableSort(PEChain_8_io_enableSort),
    .io_state(PEChain_8_io_state),
    .io_leftNBR_data(PEChain_8_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_8_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_8_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_8_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_8_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_8_io_rightNBR_compRes),
    .io_currCell_data(PEChain_8_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_8_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_8_io_currCell_compRes),
    .io_lisSize(PEChain_8_io_lisSize),
    .io_lastCell(PEChain_8_io_lastCell),
    .io_active(PEChain_8_io_active),
    .io_inData(PEChain_8_io_inData),
    .io_rightPropDiscard(PEChain_8_io_rightPropDiscard),
    .io_leftOutData(PEChain_8_io_leftOutData),
    .io_rightOutData(PEChain_8_io_rightOutData),
    .io_currDiscard(PEChain_8_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_8_io_toLeftPropDiscard)
  );
  PE_9 PEChain_9 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_9_clock),
    .reset(PEChain_9_reset),
    .io_enableSort(PEChain_9_io_enableSort),
    .io_state(PEChain_9_io_state),
    .io_leftNBR_data(PEChain_9_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_9_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_9_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_9_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_9_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_9_io_rightNBR_compRes),
    .io_currCell_data(PEChain_9_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_9_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_9_io_currCell_compRes),
    .io_lisSize(PEChain_9_io_lisSize),
    .io_lastCell(PEChain_9_io_lastCell),
    .io_active(PEChain_9_io_active),
    .io_inData(PEChain_9_io_inData),
    .io_rightPropDiscard(PEChain_9_io_rightPropDiscard),
    .io_leftOutData(PEChain_9_io_leftOutData),
    .io_rightOutData(PEChain_9_io_rightOutData),
    .io_currDiscard(PEChain_9_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_9_io_toLeftPropDiscard)
  );
  PE_10 PEChain_10 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_10_clock),
    .reset(PEChain_10_reset),
    .io_enableSort(PEChain_10_io_enableSort),
    .io_state(PEChain_10_io_state),
    .io_leftNBR_data(PEChain_10_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_10_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_10_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_10_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_10_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_10_io_rightNBR_compRes),
    .io_currCell_data(PEChain_10_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_10_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_10_io_currCell_compRes),
    .io_lisSize(PEChain_10_io_lisSize),
    .io_lastCell(PEChain_10_io_lastCell),
    .io_active(PEChain_10_io_active),
    .io_inData(PEChain_10_io_inData),
    .io_rightPropDiscard(PEChain_10_io_rightPropDiscard),
    .io_leftOutData(PEChain_10_io_leftOutData),
    .io_rightOutData(PEChain_10_io_rightOutData),
    .io_currDiscard(PEChain_10_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_10_io_toLeftPropDiscard)
  );
  PE_11 PEChain_11 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_11_clock),
    .reset(PEChain_11_reset),
    .io_enableSort(PEChain_11_io_enableSort),
    .io_state(PEChain_11_io_state),
    .io_leftNBR_data(PEChain_11_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_11_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_11_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_11_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_11_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_11_io_rightNBR_compRes),
    .io_currCell_data(PEChain_11_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_11_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_11_io_currCell_compRes),
    .io_lisSize(PEChain_11_io_lisSize),
    .io_lastCell(PEChain_11_io_lastCell),
    .io_active(PEChain_11_io_active),
    .io_inData(PEChain_11_io_inData),
    .io_rightPropDiscard(PEChain_11_io_rightPropDiscard),
    .io_leftOutData(PEChain_11_io_leftOutData),
    .io_rightOutData(PEChain_11_io_rightOutData),
    .io_currDiscard(PEChain_11_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_11_io_toLeftPropDiscard)
  );
  PE_12 PEChain_12 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_12_clock),
    .reset(PEChain_12_reset),
    .io_enableSort(PEChain_12_io_enableSort),
    .io_state(PEChain_12_io_state),
    .io_leftNBR_data(PEChain_12_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_12_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_12_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_12_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_12_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_12_io_rightNBR_compRes),
    .io_currCell_data(PEChain_12_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_12_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_12_io_currCell_compRes),
    .io_lisSize(PEChain_12_io_lisSize),
    .io_lastCell(PEChain_12_io_lastCell),
    .io_active(PEChain_12_io_active),
    .io_inData(PEChain_12_io_inData),
    .io_rightPropDiscard(PEChain_12_io_rightPropDiscard),
    .io_leftOutData(PEChain_12_io_leftOutData),
    .io_rightOutData(PEChain_12_io_rightOutData),
    .io_currDiscard(PEChain_12_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_12_io_toLeftPropDiscard)
  );
  PE_13 PEChain_13 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_13_clock),
    .reset(PEChain_13_reset),
    .io_enableSort(PEChain_13_io_enableSort),
    .io_state(PEChain_13_io_state),
    .io_leftNBR_data(PEChain_13_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_13_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_13_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_13_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_13_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_13_io_rightNBR_compRes),
    .io_currCell_data(PEChain_13_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_13_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_13_io_currCell_compRes),
    .io_lisSize(PEChain_13_io_lisSize),
    .io_lastCell(PEChain_13_io_lastCell),
    .io_active(PEChain_13_io_active),
    .io_inData(PEChain_13_io_inData),
    .io_rightPropDiscard(PEChain_13_io_rightPropDiscard),
    .io_leftOutData(PEChain_13_io_leftOutData),
    .io_rightOutData(PEChain_13_io_rightOutData),
    .io_currDiscard(PEChain_13_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_13_io_toLeftPropDiscard)
  );
  PE_14 PEChain_14 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_14_clock),
    .reset(PEChain_14_reset),
    .io_enableSort(PEChain_14_io_enableSort),
    .io_state(PEChain_14_io_state),
    .io_leftNBR_data(PEChain_14_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_14_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_14_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_14_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_14_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_14_io_rightNBR_compRes),
    .io_currCell_data(PEChain_14_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_14_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_14_io_currCell_compRes),
    .io_lisSize(PEChain_14_io_lisSize),
    .io_lastCell(PEChain_14_io_lastCell),
    .io_active(PEChain_14_io_active),
    .io_inData(PEChain_14_io_inData),
    .io_rightPropDiscard(PEChain_14_io_rightPropDiscard),
    .io_leftOutData(PEChain_14_io_leftOutData),
    .io_rightOutData(PEChain_14_io_rightOutData),
    .io_currDiscard(PEChain_14_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_14_io_toLeftPropDiscard)
  );
  PE_15 PEChain_15 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_15_clock),
    .reset(PEChain_15_reset),
    .io_enableSort(PEChain_15_io_enableSort),
    .io_state(PEChain_15_io_state),
    .io_leftNBR_data(PEChain_15_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_15_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_15_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_15_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_15_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_15_io_rightNBR_compRes),
    .io_currCell_data(PEChain_15_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_15_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_15_io_currCell_compRes),
    .io_lisSize(PEChain_15_io_lisSize),
    .io_lastCell(PEChain_15_io_lastCell),
    .io_active(PEChain_15_io_active),
    .io_inData(PEChain_15_io_inData),
    .io_rightPropDiscard(PEChain_15_io_rightPropDiscard),
    .io_leftOutData(PEChain_15_io_leftOutData),
    .io_rightOutData(PEChain_15_io_rightOutData),
    .io_currDiscard(PEChain_15_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_15_io_toLeftPropDiscard)
  );
  PE_16 PEChain_16 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_16_clock),
    .reset(PEChain_16_reset),
    .io_enableSort(PEChain_16_io_enableSort),
    .io_state(PEChain_16_io_state),
    .io_leftNBR_data(PEChain_16_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_16_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_16_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_16_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_16_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_16_io_rightNBR_compRes),
    .io_currCell_data(PEChain_16_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_16_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_16_io_currCell_compRes),
    .io_lisSize(PEChain_16_io_lisSize),
    .io_lastCell(PEChain_16_io_lastCell),
    .io_active(PEChain_16_io_active),
    .io_inData(PEChain_16_io_inData),
    .io_rightPropDiscard(PEChain_16_io_rightPropDiscard),
    .io_leftOutData(PEChain_16_io_leftOutData),
    .io_rightOutData(PEChain_16_io_rightOutData),
    .io_currDiscard(PEChain_16_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_16_io_toLeftPropDiscard)
  );
  PE_17 PEChain_17 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_17_clock),
    .reset(PEChain_17_reset),
    .io_enableSort(PEChain_17_io_enableSort),
    .io_state(PEChain_17_io_state),
    .io_leftNBR_data(PEChain_17_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_17_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_17_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_17_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_17_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_17_io_rightNBR_compRes),
    .io_currCell_data(PEChain_17_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_17_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_17_io_currCell_compRes),
    .io_lisSize(PEChain_17_io_lisSize),
    .io_lastCell(PEChain_17_io_lastCell),
    .io_active(PEChain_17_io_active),
    .io_inData(PEChain_17_io_inData),
    .io_rightPropDiscard(PEChain_17_io_rightPropDiscard),
    .io_leftOutData(PEChain_17_io_leftOutData),
    .io_rightOutData(PEChain_17_io_rightOutData),
    .io_currDiscard(PEChain_17_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_17_io_toLeftPropDiscard)
  );
  PE_18 PEChain_18 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_18_clock),
    .reset(PEChain_18_reset),
    .io_enableSort(PEChain_18_io_enableSort),
    .io_state(PEChain_18_io_state),
    .io_leftNBR_data(PEChain_18_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_18_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_18_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_18_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_18_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_18_io_rightNBR_compRes),
    .io_currCell_data(PEChain_18_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_18_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_18_io_currCell_compRes),
    .io_lisSize(PEChain_18_io_lisSize),
    .io_lastCell(PEChain_18_io_lastCell),
    .io_active(PEChain_18_io_active),
    .io_inData(PEChain_18_io_inData),
    .io_rightPropDiscard(PEChain_18_io_rightPropDiscard),
    .io_leftOutData(PEChain_18_io_leftOutData),
    .io_rightOutData(PEChain_18_io_rightOutData),
    .io_currDiscard(PEChain_18_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_18_io_toLeftPropDiscard)
  );
  PE_19 PEChain_19 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_19_clock),
    .reset(PEChain_19_reset),
    .io_enableSort(PEChain_19_io_enableSort),
    .io_state(PEChain_19_io_state),
    .io_leftNBR_data(PEChain_19_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_19_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_19_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_19_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_19_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_19_io_rightNBR_compRes),
    .io_currCell_data(PEChain_19_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_19_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_19_io_currCell_compRes),
    .io_lisSize(PEChain_19_io_lisSize),
    .io_lastCell(PEChain_19_io_lastCell),
    .io_active(PEChain_19_io_active),
    .io_inData(PEChain_19_io_inData),
    .io_rightPropDiscard(PEChain_19_io_rightPropDiscard),
    .io_leftOutData(PEChain_19_io_leftOutData),
    .io_rightOutData(PEChain_19_io_rightOutData),
    .io_currDiscard(PEChain_19_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_19_io_toLeftPropDiscard)
  );
  PE_20 PEChain_20 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_20_clock),
    .reset(PEChain_20_reset),
    .io_enableSort(PEChain_20_io_enableSort),
    .io_state(PEChain_20_io_state),
    .io_leftNBR_data(PEChain_20_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_20_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_20_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_20_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_20_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_20_io_rightNBR_compRes),
    .io_currCell_data(PEChain_20_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_20_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_20_io_currCell_compRes),
    .io_lisSize(PEChain_20_io_lisSize),
    .io_lastCell(PEChain_20_io_lastCell),
    .io_active(PEChain_20_io_active),
    .io_inData(PEChain_20_io_inData),
    .io_rightPropDiscard(PEChain_20_io_rightPropDiscard),
    .io_leftOutData(PEChain_20_io_leftOutData),
    .io_rightOutData(PEChain_20_io_rightOutData),
    .io_currDiscard(PEChain_20_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_20_io_toLeftPropDiscard)
  );
  PE_21 PEChain_21 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_21_clock),
    .reset(PEChain_21_reset),
    .io_enableSort(PEChain_21_io_enableSort),
    .io_state(PEChain_21_io_state),
    .io_leftNBR_data(PEChain_21_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_21_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_21_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_21_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_21_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_21_io_rightNBR_compRes),
    .io_currCell_data(PEChain_21_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_21_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_21_io_currCell_compRes),
    .io_lisSize(PEChain_21_io_lisSize),
    .io_lastCell(PEChain_21_io_lastCell),
    .io_active(PEChain_21_io_active),
    .io_inData(PEChain_21_io_inData),
    .io_rightPropDiscard(PEChain_21_io_rightPropDiscard),
    .io_leftOutData(PEChain_21_io_leftOutData),
    .io_rightOutData(PEChain_21_io_rightOutData),
    .io_currDiscard(PEChain_21_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_21_io_toLeftPropDiscard)
  );
  PE_22 PEChain_22 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_22_clock),
    .reset(PEChain_22_reset),
    .io_enableSort(PEChain_22_io_enableSort),
    .io_state(PEChain_22_io_state),
    .io_leftNBR_data(PEChain_22_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_22_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_22_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_22_io_rightNBR_data),
    .io_rightNBR_lifeCNT(PEChain_22_io_rightNBR_lifeCNT),
    .io_rightNBR_compRes(PEChain_22_io_rightNBR_compRes),
    .io_currCell_data(PEChain_22_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_22_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_22_io_currCell_compRes),
    .io_lisSize(PEChain_22_io_lisSize),
    .io_lastCell(PEChain_22_io_lastCell),
    .io_active(PEChain_22_io_active),
    .io_inData(PEChain_22_io_inData),
    .io_rightPropDiscard(PEChain_22_io_rightPropDiscard),
    .io_leftOutData(PEChain_22_io_leftOutData),
    .io_rightOutData(PEChain_22_io_rightOutData),
    .io_currDiscard(PEChain_22_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_22_io_toLeftPropDiscard)
  );
  PE_23 PEChain_23 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_23_clock),
    .reset(PEChain_23_reset),
    .io_enableSort(PEChain_23_io_enableSort),
    .io_state(PEChain_23_io_state),
    .io_leftNBR_data(PEChain_23_io_leftNBR_data),
    .io_leftNBR_lifeCNT(PEChain_23_io_leftNBR_lifeCNT),
    .io_leftNBR_compRes(PEChain_23_io_leftNBR_compRes),
    .io_currCell_data(PEChain_23_io_currCell_data),
    .io_currCell_lifeCNT(PEChain_23_io_currCell_lifeCNT),
    .io_currCell_compRes(PEChain_23_io_currCell_compRes),
    .io_lisSize(PEChain_23_io_lisSize),
    .io_lastCell(PEChain_23_io_lastCell),
    .io_active(PEChain_23_io_active),
    .io_inData(PEChain_23_io_inData),
    .io_leftOutData(PEChain_23_io_leftOutData),
    .io_currDiscard(PEChain_23_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_23_io_toLeftPropDiscard)
  );
  assign _T_1 = lisSizeReg - 6'h1; // @[LinearSorter.scala 86:43]
  assign _T_96 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_98 = cntInData + 5'h1; // @[LinearSorter.scala 92:28]
  assign _T_99 = state == 2'h0; // @[LinearSorter.scala 94:20]
  assign _GEN_39 = {{1'd0}, cntInData}; // @[LinearSorter.scala 98:19]
  assign _T_102 = _GEN_39 == _T_1; // @[LinearSorter.scala 98:19]
  assign _T_104 = _T_102 & _T_96; // @[LinearSorter.scala 98:42]
  assign _T_113 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_7 = _T_96 ? 2'h1 : state; // @[LinearSorter.scala 117:27]
  assign _T_115 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign fireLastIn = io_lastIn & _T_96; // @[LinearSorter.scala 111:30]
  assign _GEN_8 = fireLastIn ? 2'h2 : state; // @[LinearSorter.scala 120:62]
  assign _T_117 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_40 = {{1'd0}, cntOutData}; // @[LinearSorter.scala 125:28]
  assign _T_120 = _GEN_40 == _T_1; // @[LinearSorter.scala 125:28]
  assign _GEN_9 = _T_120 ? 2'h0 : state; // @[LinearSorter.scala 125:50]
  assign _GEN_10 = _T_117 ? _GEN_9 : state; // @[Conditional.scala 39:67]
  assign _GEN_11 = _T_115 ? _GEN_8 : _GEN_10; // @[Conditional.scala 39:67]
  assign state_next = _T_113 ? _GEN_7 : _GEN_11; // @[Conditional.scala 40:58]
  assign _T_105 = state_next == 2'h0; // @[LinearSorter.scala 101:25]
  assign _GEN_2 = _T_105 ? 1'h0 : initialInDone; // @[LinearSorter.scala 101:36]
  assign _GEN_3 = _T_104 | _GEN_2; // @[LinearSorter.scala 98:59]
  assign _T_106 = io_out_valid & io_out_ready; // @[LinearSorter.scala 106:29]
  assign _T_107 = state == 2'h2; // @[LinearSorter.scala 106:54]
  assign enable = _T_106 & _T_107; // @[LinearSorter.scala 106:45]
  assign _T_109 = cntOutData == 5'h17; // @[LISutil.scala 13:24]
  assign _T_111 = cntOutData + 5'h1; // @[LISutil.scala 14:22]
  assign _T_126 = _T_107 & io_out_ready; // @[LinearSorter.scala 168:63]
  assign discardSignals_2 = PEChain_2_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_1 = PEChain_1_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_0 = PEChain_0_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_5 = PEChain_5_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_4 = PEChain_4_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_3 = PEChain_3_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_293 = {discardSignals_5,discardSignals_4,discardSignals_3,discardSignals_2,discardSignals_1,discardSignals_0}; // @[LinearSorter.scala 177:50]
  assign discardSignals_8 = PEChain_8_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_7 = PEChain_7_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_6 = PEChain_6_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_11 = PEChain_11_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_10 = PEChain_10_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_9 = PEChain_9_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_299 = {discardSignals_11,discardSignals_10,discardSignals_9,discardSignals_8,discardSignals_7,discardSignals_6,_T_293}; // @[LinearSorter.scala 177:50]
  assign discardSignals_14 = PEChain_14_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_13 = PEChain_13_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_12 = PEChain_12_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_17 = PEChain_17_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_16 = PEChain_16_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_15 = PEChain_15_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_304 = {discardSignals_17,discardSignals_16,discardSignals_15,discardSignals_14,discardSignals_13,discardSignals_12}; // @[LinearSorter.scala 177:50]
  assign discardSignals_20 = PEChain_20_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_19 = PEChain_19_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_18 = PEChain_18_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_23 = PEChain_23_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_22 = PEChain_22_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_21 = PEChain_21_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_311 = {discardSignals_23,discardSignals_22,discardSignals_21,discardSignals_20,discardSignals_19,discardSignals_18,_T_304,_T_299}; // @[LinearSorter.scala 177:50]
  assign _T_336 = _T_311[22] ? 5'h16 : 5'h17; // @[Mux.scala 47:69]
  assign _T_337 = _T_311[21] ? 5'h15 : _T_336; // @[Mux.scala 47:69]
  assign _T_338 = _T_311[20] ? 5'h14 : _T_337; // @[Mux.scala 47:69]
  assign _T_339 = _T_311[19] ? 5'h13 : _T_338; // @[Mux.scala 47:69]
  assign _T_340 = _T_311[18] ? 5'h12 : _T_339; // @[Mux.scala 47:69]
  assign _T_341 = _T_311[17] ? 5'h11 : _T_340; // @[Mux.scala 47:69]
  assign _T_342 = _T_311[16] ? 5'h10 : _T_341; // @[Mux.scala 47:69]
  assign _T_343 = _T_311[15] ? 5'hf : _T_342; // @[Mux.scala 47:69]
  assign _T_344 = _T_311[14] ? 5'he : _T_343; // @[Mux.scala 47:69]
  assign _T_345 = _T_311[13] ? 5'hd : _T_344; // @[Mux.scala 47:69]
  assign _T_346 = _T_311[12] ? 5'hc : _T_345; // @[Mux.scala 47:69]
  assign _T_347 = _T_311[11] ? 5'hb : _T_346; // @[Mux.scala 47:69]
  assign _T_348 = _T_311[10] ? 5'ha : _T_347; // @[Mux.scala 47:69]
  assign _T_349 = _T_311[9] ? 5'h9 : _T_348; // @[Mux.scala 47:69]
  assign _T_350 = _T_311[8] ? 5'h8 : _T_349; // @[Mux.scala 47:69]
  assign _T_351 = _T_311[7] ? 5'h7 : _T_350; // @[Mux.scala 47:69]
  assign _T_352 = _T_311[6] ? 5'h6 : _T_351; // @[Mux.scala 47:69]
  assign _T_353 = _T_311[5] ? 5'h5 : _T_352; // @[Mux.scala 47:69]
  assign _T_354 = _T_311[4] ? 5'h4 : _T_353; // @[Mux.scala 47:69]
  assign _T_355 = _T_311[3] ? 5'h3 : _T_354; // @[Mux.scala 47:69]
  assign _T_356 = _T_311[2] ? 5'h2 : _T_355; // @[Mux.scala 47:69]
  assign _T_357 = _T_311[1] ? 5'h1 : _T_356; // @[Mux.scala 47:69]
  assign getDiscarded = _T_311[0] ? 5'h0 : _T_357; // @[Mux.scala 47:69]
  assign _T_359 = state != 2'h2; // @[LinearSorter.scala 199:49]
  assign outputData_0 = PEChain_0_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign outputData_1 = PEChain_1_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_16 = 5'h1 == getDiscarded ? $signed(outputData_1) : $signed(outputData_0); // @[LinearSorter.scala 206:15]
  assign outputData_2 = PEChain_2_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_17 = 5'h2 == getDiscarded ? $signed(outputData_2) : $signed(_GEN_16); // @[LinearSorter.scala 206:15]
  assign outputData_3 = PEChain_3_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_18 = 5'h3 == getDiscarded ? $signed(outputData_3) : $signed(_GEN_17); // @[LinearSorter.scala 206:15]
  assign outputData_4 = PEChain_4_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_19 = 5'h4 == getDiscarded ? $signed(outputData_4) : $signed(_GEN_18); // @[LinearSorter.scala 206:15]
  assign outputData_5 = PEChain_5_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_20 = 5'h5 == getDiscarded ? $signed(outputData_5) : $signed(_GEN_19); // @[LinearSorter.scala 206:15]
  assign outputData_6 = PEChain_6_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_21 = 5'h6 == getDiscarded ? $signed(outputData_6) : $signed(_GEN_20); // @[LinearSorter.scala 206:15]
  assign outputData_7 = PEChain_7_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_22 = 5'h7 == getDiscarded ? $signed(outputData_7) : $signed(_GEN_21); // @[LinearSorter.scala 206:15]
  assign outputData_8 = PEChain_8_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_23 = 5'h8 == getDiscarded ? $signed(outputData_8) : $signed(_GEN_22); // @[LinearSorter.scala 206:15]
  assign outputData_9 = PEChain_9_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_24 = 5'h9 == getDiscarded ? $signed(outputData_9) : $signed(_GEN_23); // @[LinearSorter.scala 206:15]
  assign outputData_10 = PEChain_10_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_25 = 5'ha == getDiscarded ? $signed(outputData_10) : $signed(_GEN_24); // @[LinearSorter.scala 206:15]
  assign outputData_11 = PEChain_11_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_26 = 5'hb == getDiscarded ? $signed(outputData_11) : $signed(_GEN_25); // @[LinearSorter.scala 206:15]
  assign outputData_12 = PEChain_12_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_27 = 5'hc == getDiscarded ? $signed(outputData_12) : $signed(_GEN_26); // @[LinearSorter.scala 206:15]
  assign outputData_13 = PEChain_13_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_28 = 5'hd == getDiscarded ? $signed(outputData_13) : $signed(_GEN_27); // @[LinearSorter.scala 206:15]
  assign outputData_14 = PEChain_14_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_29 = 5'he == getDiscarded ? $signed(outputData_14) : $signed(_GEN_28); // @[LinearSorter.scala 206:15]
  assign outputData_15 = PEChain_15_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_30 = 5'hf == getDiscarded ? $signed(outputData_15) : $signed(_GEN_29); // @[LinearSorter.scala 206:15]
  assign outputData_16 = PEChain_16_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_31 = 5'h10 == getDiscarded ? $signed(outputData_16) : $signed(_GEN_30); // @[LinearSorter.scala 206:15]
  assign outputData_17 = PEChain_17_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_32 = 5'h11 == getDiscarded ? $signed(outputData_17) : $signed(_GEN_31); // @[LinearSorter.scala 206:15]
  assign outputData_18 = PEChain_18_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_33 = 5'h12 == getDiscarded ? $signed(outputData_18) : $signed(_GEN_32); // @[LinearSorter.scala 206:15]
  assign outputData_19 = PEChain_19_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_34 = 5'h13 == getDiscarded ? $signed(outputData_19) : $signed(_GEN_33); // @[LinearSorter.scala 206:15]
  assign outputData_20 = PEChain_20_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_35 = 5'h14 == getDiscarded ? $signed(outputData_20) : $signed(_GEN_34); // @[LinearSorter.scala 206:15]
  assign outputData_21 = PEChain_21_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_36 = 5'h15 == getDiscarded ? $signed(outputData_21) : $signed(_GEN_35); // @[LinearSorter.scala 206:15]
  assign outputData_22 = PEChain_22_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_37 = 5'h16 == getDiscarded ? $signed(outputData_22) : $signed(_GEN_36); // @[LinearSorter.scala 206:15]
  assign outputData_23 = PEChain_23_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _T_365 = ~initialInDone; // @[LinearSorter.scala 208:18]
  assign _T_367 = io_out_ready & _T_359; // @[LinearSorter.scala 208:49]
  assign _T_369 = initialInDone & io_in_valid; // @[LinearSorter.scala 209:33]
  assign io_in_ready = _T_365 | _T_367; // @[LinearSorter.scala 208:15]
  assign io_out_valid = _T_369 | _T_107; // @[LinearSorter.scala 209:16]
  assign io_out_bits = 5'h17 == getDiscarded ? $signed(outputData_23) : $signed(_GEN_37); // @[LinearSorter.scala 206:15]
  assign io_lastOut = _GEN_40 == _T_1; // @[LinearSorter.scala 207:15]
  assign io_sortedData_0 = PEChain_0_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_1 = PEChain_1_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_2 = PEChain_2_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_3 = PEChain_3_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_4 = PEChain_4_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_5 = PEChain_5_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_6 = PEChain_6_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_7 = PEChain_7_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_8 = PEChain_8_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_9 = PEChain_9_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_10 = PEChain_10_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_11 = PEChain_11_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_12 = PEChain_12_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_13 = PEChain_13_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_14 = PEChain_14_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_15 = PEChain_15_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_16 = PEChain_16_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_17 = PEChain_17_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_18 = PEChain_18_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_19 = PEChain_19_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_20 = PEChain_20_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_21 = PEChain_21_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_22 = PEChain_22_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_23 = PEChain_23_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sorterFull = initialInDone & _T_359; // @[LinearSorter.scala 199:23]
  assign io_sorterEmpty = state == 2'h0; // @[LinearSorter.scala 202:24]
  assign PEChain_0_clock = clock;
  assign PEChain_0_reset = reset;
  assign PEChain_0_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_0_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_0_io_rightNBR_data = PEChain_1_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_0_io_rightNBR_lifeCNT = PEChain_1_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_0_io_rightNBR_compRes = PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_0_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_0_io_lastCell = 6'h0 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_0_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_0_io_rightPropDiscard = PEChain_1_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_1_clock = clock;
  assign PEChain_1_reset = reset;
  assign PEChain_1_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_1_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_1_io_leftNBR_data = PEChain_0_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_1_io_leftNBR_lifeCNT = PEChain_0_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_1_io_leftNBR_compRes = PEChain_0_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_1_io_rightNBR_data = PEChain_2_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_1_io_rightNBR_lifeCNT = PEChain_2_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_1_io_rightNBR_compRes = PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_1_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_1_io_lastCell = 6'h1 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_1_io_active = 6'h1 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_1_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_1_io_rightPropDiscard = PEChain_2_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_2_clock = clock;
  assign PEChain_2_reset = reset;
  assign PEChain_2_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_2_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_2_io_leftNBR_data = PEChain_1_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_2_io_leftNBR_lifeCNT = PEChain_1_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_2_io_leftNBR_compRes = PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_2_io_rightNBR_data = PEChain_3_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_2_io_rightNBR_lifeCNT = PEChain_3_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_2_io_rightNBR_compRes = PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_2_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_2_io_lastCell = 6'h2 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_2_io_active = 6'h2 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_2_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_2_io_rightPropDiscard = PEChain_3_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_3_clock = clock;
  assign PEChain_3_reset = reset;
  assign PEChain_3_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_3_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_3_io_leftNBR_data = PEChain_2_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_3_io_leftNBR_lifeCNT = PEChain_2_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_3_io_leftNBR_compRes = PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_3_io_rightNBR_data = PEChain_4_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_3_io_rightNBR_lifeCNT = PEChain_4_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_3_io_rightNBR_compRes = PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_3_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_3_io_lastCell = 6'h3 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_3_io_active = 6'h3 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_3_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_3_io_rightPropDiscard = PEChain_4_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_4_clock = clock;
  assign PEChain_4_reset = reset;
  assign PEChain_4_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_4_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_4_io_leftNBR_data = PEChain_3_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_4_io_leftNBR_lifeCNT = PEChain_3_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_4_io_leftNBR_compRes = PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_4_io_rightNBR_data = PEChain_5_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_4_io_rightNBR_lifeCNT = PEChain_5_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_4_io_rightNBR_compRes = PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_4_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_4_io_lastCell = 6'h4 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_4_io_active = 6'h4 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_4_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_4_io_rightPropDiscard = PEChain_5_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_5_clock = clock;
  assign PEChain_5_reset = reset;
  assign PEChain_5_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_5_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_5_io_leftNBR_data = PEChain_4_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_5_io_leftNBR_lifeCNT = PEChain_4_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_5_io_leftNBR_compRes = PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_5_io_rightNBR_data = PEChain_6_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_5_io_rightNBR_lifeCNT = PEChain_6_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_5_io_rightNBR_compRes = PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_5_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_5_io_lastCell = 6'h5 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_5_io_active = 6'h5 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_5_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_5_io_rightPropDiscard = PEChain_6_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_6_clock = clock;
  assign PEChain_6_reset = reset;
  assign PEChain_6_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_6_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_6_io_leftNBR_data = PEChain_5_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_6_io_leftNBR_lifeCNT = PEChain_5_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_6_io_leftNBR_compRes = PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_6_io_rightNBR_data = PEChain_7_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_6_io_rightNBR_lifeCNT = PEChain_7_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_6_io_rightNBR_compRes = PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_6_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_6_io_lastCell = 6'h6 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_6_io_active = 6'h6 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_6_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_6_io_rightPropDiscard = PEChain_7_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_7_clock = clock;
  assign PEChain_7_reset = reset;
  assign PEChain_7_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_7_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_7_io_leftNBR_data = PEChain_6_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_7_io_leftNBR_lifeCNT = PEChain_6_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_7_io_leftNBR_compRes = PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_7_io_rightNBR_data = PEChain_8_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_7_io_rightNBR_lifeCNT = PEChain_8_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_7_io_rightNBR_compRes = PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_7_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_7_io_lastCell = 6'h7 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_7_io_active = 6'h7 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_7_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_7_io_rightPropDiscard = PEChain_8_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_8_clock = clock;
  assign PEChain_8_reset = reset;
  assign PEChain_8_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_8_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_8_io_leftNBR_data = PEChain_7_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_8_io_leftNBR_lifeCNT = PEChain_7_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_8_io_leftNBR_compRes = PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_8_io_rightNBR_data = PEChain_9_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_8_io_rightNBR_lifeCNT = PEChain_9_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_8_io_rightNBR_compRes = PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_8_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_8_io_lastCell = 6'h8 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_8_io_active = 6'h8 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_8_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_8_io_rightPropDiscard = PEChain_9_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_9_clock = clock;
  assign PEChain_9_reset = reset;
  assign PEChain_9_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_9_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_9_io_leftNBR_data = PEChain_8_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_9_io_leftNBR_lifeCNT = PEChain_8_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_9_io_leftNBR_compRes = PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_9_io_rightNBR_data = PEChain_10_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_9_io_rightNBR_lifeCNT = PEChain_10_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_9_io_rightNBR_compRes = PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_9_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_9_io_lastCell = 6'h9 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_9_io_active = 6'h9 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_9_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_9_io_rightPropDiscard = PEChain_10_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_10_clock = clock;
  assign PEChain_10_reset = reset;
  assign PEChain_10_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_10_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_10_io_leftNBR_data = PEChain_9_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_10_io_leftNBR_lifeCNT = PEChain_9_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_10_io_leftNBR_compRes = PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_10_io_rightNBR_data = PEChain_11_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_10_io_rightNBR_lifeCNT = PEChain_11_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_10_io_rightNBR_compRes = PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_10_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_10_io_lastCell = 6'ha == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_10_io_active = 6'ha <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_10_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_10_io_rightPropDiscard = PEChain_11_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_11_clock = clock;
  assign PEChain_11_reset = reset;
  assign PEChain_11_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_11_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_11_io_leftNBR_data = PEChain_10_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_11_io_leftNBR_lifeCNT = PEChain_10_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_11_io_leftNBR_compRes = PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_11_io_rightNBR_data = PEChain_12_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_11_io_rightNBR_lifeCNT = PEChain_12_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_11_io_rightNBR_compRes = PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_11_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_11_io_lastCell = 6'hb == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_11_io_active = 6'hb <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_11_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_11_io_rightPropDiscard = PEChain_12_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_12_clock = clock;
  assign PEChain_12_reset = reset;
  assign PEChain_12_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_12_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_12_io_leftNBR_data = PEChain_11_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_12_io_leftNBR_lifeCNT = PEChain_11_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_12_io_leftNBR_compRes = PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_12_io_rightNBR_data = PEChain_13_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_12_io_rightNBR_lifeCNT = PEChain_13_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_12_io_rightNBR_compRes = PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_12_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_12_io_lastCell = 6'hc == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_12_io_active = 6'hc <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_12_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_12_io_rightPropDiscard = PEChain_13_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_13_clock = clock;
  assign PEChain_13_reset = reset;
  assign PEChain_13_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_13_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_13_io_leftNBR_data = PEChain_12_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_13_io_leftNBR_lifeCNT = PEChain_12_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_13_io_leftNBR_compRes = PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_13_io_rightNBR_data = PEChain_14_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_13_io_rightNBR_lifeCNT = PEChain_14_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_13_io_rightNBR_compRes = PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_13_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_13_io_lastCell = 6'hd == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_13_io_active = 6'hd <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_13_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_13_io_rightPropDiscard = PEChain_14_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_14_clock = clock;
  assign PEChain_14_reset = reset;
  assign PEChain_14_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_14_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_14_io_leftNBR_data = PEChain_13_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_14_io_leftNBR_lifeCNT = PEChain_13_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_14_io_leftNBR_compRes = PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_14_io_rightNBR_data = PEChain_15_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_14_io_rightNBR_lifeCNT = PEChain_15_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_14_io_rightNBR_compRes = PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_14_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_14_io_lastCell = 6'he == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_14_io_active = 6'he <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_14_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_14_io_rightPropDiscard = PEChain_15_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_15_clock = clock;
  assign PEChain_15_reset = reset;
  assign PEChain_15_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_15_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_15_io_leftNBR_data = PEChain_14_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_15_io_leftNBR_lifeCNT = PEChain_14_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_15_io_leftNBR_compRes = PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_15_io_rightNBR_data = PEChain_16_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_15_io_rightNBR_lifeCNT = PEChain_16_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_15_io_rightNBR_compRes = PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_15_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_15_io_lastCell = 6'hf == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_15_io_active = 6'hf <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_15_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_15_io_rightPropDiscard = PEChain_16_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_16_clock = clock;
  assign PEChain_16_reset = reset;
  assign PEChain_16_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_16_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_16_io_leftNBR_data = PEChain_15_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_16_io_leftNBR_lifeCNT = PEChain_15_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_16_io_leftNBR_compRes = PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_16_io_rightNBR_data = PEChain_17_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_16_io_rightNBR_lifeCNT = PEChain_17_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_16_io_rightNBR_compRes = PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_16_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_16_io_lastCell = 6'h10 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_16_io_active = 6'h10 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_16_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_16_io_rightPropDiscard = PEChain_17_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_17_clock = clock;
  assign PEChain_17_reset = reset;
  assign PEChain_17_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_17_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_17_io_leftNBR_data = PEChain_16_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_17_io_leftNBR_lifeCNT = PEChain_16_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_17_io_leftNBR_compRes = PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_17_io_rightNBR_data = PEChain_18_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_17_io_rightNBR_lifeCNT = PEChain_18_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_17_io_rightNBR_compRes = PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_17_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_17_io_lastCell = 6'h11 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_17_io_active = 6'h11 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_17_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_17_io_rightPropDiscard = PEChain_18_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_18_clock = clock;
  assign PEChain_18_reset = reset;
  assign PEChain_18_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_18_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_18_io_leftNBR_data = PEChain_17_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_18_io_leftNBR_lifeCNT = PEChain_17_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_18_io_leftNBR_compRes = PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_18_io_rightNBR_data = PEChain_19_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_18_io_rightNBR_lifeCNT = PEChain_19_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_18_io_rightNBR_compRes = PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_18_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_18_io_lastCell = 6'h12 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_18_io_active = 6'h12 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_18_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_18_io_rightPropDiscard = PEChain_19_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_19_clock = clock;
  assign PEChain_19_reset = reset;
  assign PEChain_19_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_19_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_19_io_leftNBR_data = PEChain_18_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_19_io_leftNBR_lifeCNT = PEChain_18_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_19_io_leftNBR_compRes = PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_19_io_rightNBR_data = PEChain_20_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_19_io_rightNBR_lifeCNT = PEChain_20_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_19_io_rightNBR_compRes = PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_19_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_19_io_lastCell = 6'h13 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_19_io_active = 6'h13 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_19_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_19_io_rightPropDiscard = PEChain_20_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_20_clock = clock;
  assign PEChain_20_reset = reset;
  assign PEChain_20_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_20_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_20_io_leftNBR_data = PEChain_19_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_20_io_leftNBR_lifeCNT = PEChain_19_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_20_io_leftNBR_compRes = PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_20_io_rightNBR_data = PEChain_21_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_20_io_rightNBR_lifeCNT = PEChain_21_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_20_io_rightNBR_compRes = PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_20_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_20_io_lastCell = 6'h14 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_20_io_active = 6'h14 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_20_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_20_io_rightPropDiscard = PEChain_21_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_21_clock = clock;
  assign PEChain_21_reset = reset;
  assign PEChain_21_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_21_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_21_io_leftNBR_data = PEChain_20_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_21_io_leftNBR_lifeCNT = PEChain_20_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_21_io_leftNBR_compRes = PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_21_io_rightNBR_data = PEChain_22_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_21_io_rightNBR_lifeCNT = PEChain_22_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_21_io_rightNBR_compRes = PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_21_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_21_io_lastCell = 6'h15 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_21_io_active = 6'h15 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_21_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_21_io_rightPropDiscard = PEChain_22_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_22_clock = clock;
  assign PEChain_22_reset = reset;
  assign PEChain_22_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_22_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_22_io_leftNBR_data = PEChain_21_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_22_io_leftNBR_lifeCNT = PEChain_21_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_22_io_leftNBR_compRes = PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_22_io_rightNBR_data = PEChain_23_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_22_io_rightNBR_lifeCNT = PEChain_23_io_currCell_lifeCNT; // @[LinearSorter.scala 192:33]
  assign PEChain_22_io_rightNBR_compRes = PEChain_23_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_22_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_22_io_lastCell = 6'h16 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_22_io_active = 6'h16 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_22_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
  assign PEChain_22_io_rightPropDiscard = PEChain_23_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_23_clock = clock;
  assign PEChain_23_reset = reset;
  assign PEChain_23_io_enableSort = _T_96 | _T_126; // @[LinearSorter.scala 168:26]
  assign PEChain_23_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_23_io_leftNBR_data = PEChain_22_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_23_io_leftNBR_lifeCNT = PEChain_22_io_currCell_lifeCNT; // @[LinearSorter.scala 189:32]
  assign PEChain_23_io_leftNBR_compRes = PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_23_io_lisSize = io_lisSize; // @[LinearSorter.scala 146:29]
  assign PEChain_23_io_lastCell = 6'h17 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_23_io_active = 6'h17 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_23_io_inData = io_in_bits; // @[LinearSorter.scala 144:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntInData = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  lisSizeReg = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cntOutData = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_3;
    end
    if (reset) begin
      cntInData <= 5'h0;
    end else if (_T_96) begin
      cntInData <= _T_98;
    end else if (_T_99) begin
      cntInData <= 5'h0;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_113) begin
      if (_T_96) begin
        state <= 2'h1;
      end
    end else if (_T_115) begin
      if (fireLastIn) begin
        state <= 2'h2;
      end
    end else if (_T_117) begin
      if (_T_120) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      lisSizeReg <= 6'h18;
    end else if (_T_113) begin
      lisSizeReg <= io_lisSize;
    end
    if (reset) begin
      cntOutData <= 5'h0;
    end else if (_T_99) begin
      cntOutData <= 5'h0;
    end else if (enable) begin
      if (_T_109) begin
        cntOutData <= 5'h0;
      end else begin
        cntOutData <= _T_111;
      end
    end
  end
endmodule
module AXI4LISBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  lis_clock; // @[LISDspBlock.scala 55:21]
  wire  lis_reset; // @[LISDspBlock.scala 55:21]
  wire  lis_io_in_ready; // @[LISDspBlock.scala 55:21]
  wire  lis_io_in_valid; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_in_bits; // @[LISDspBlock.scala 55:21]
  wire  lis_io_lastIn; // @[LISDspBlock.scala 55:21]
  wire  lis_io_out_ready; // @[LISDspBlock.scala 55:21]
  wire  lis_io_out_valid; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_out_bits; // @[LISDspBlock.scala 55:21]
  wire  lis_io_lastOut; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_0; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_1; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_2; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_3; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_4; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_5; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_6; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_7; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_8; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_9; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_10; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_11; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_12; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_13; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_14; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_15; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_16; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_17; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_18; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_19; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_20; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_21; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_22; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_23; // @[LISDspBlock.scala 55:21]
  wire  lis_io_sorterFull; // @[LISDspBlock.scala 55:21]
  wire  lis_io_sorterEmpty; // @[LISDspBlock.scala 55:21]
  wire [5:0] lis_io_lisSize; // @[LISDspBlock.scala 55:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  sortDir; // @[LISDspBlock.scala 58:26]
  reg [31:0] _RAND_0;
  reg  flushData; // @[LISDspBlock.scala 59:28]
  reg [31:0] _RAND_1;
  reg [4:0] discardPos; // @[LISDspBlock.scala 60:29]
  reg [31:0] _RAND_2;
  reg [4:0] sendOnOutput; // @[LISDspBlock.scala 61:31]
  reg [31:0] _RAND_3;
  reg [4:0] lisSize; // @[LISDspBlock.scala 62:26]
  reg [31:0] _RAND_4;
  reg  sorterFull; // @[LISDspBlock.scala 65:29]
  reg [31:0] _RAND_5;
  reg  sorterEmpty; // @[LISDspBlock.scala 66:30]
  reg [31:0] _RAND_6;
  wire [31:0] _T_2; // @[LISDspBlock.scala 71:44]
  wire [15:0] _GEN_0; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_1; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_2; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_3; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_4; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_5; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_6; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_7; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_8; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_9; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_10; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_11; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_12; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_13; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_14; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_15; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_16; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_17; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_18; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_19; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_20; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_21; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_22; // @[LISDspBlock.scala 92:82]
  wire [15:0] _T_4; // @[LISDspBlock.scala 92:82]
  wire  _T_7; // @[RegisterRouter.scala 40:39]
  wire  _T_8; // @[RegisterRouter.scala 40:26]
  wire  _T_9; // @[RegisterRouter.scala 42:29]
  wire  _T_52_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_16; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_281; // @[Cat.scala 29:58]
  wire [5:0] _T_56; // @[RegisterRouter.scala 59:16]
  wire  _T_64; // @[RegisterRouter.scala 59:16]
  wire  _T_10; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_19; // @[OneHot.scala 65:12]
  wire [1:0] _T_21; // @[Misc.scala 200:81]
  wire  _T_22; // @[Misc.scala 204:21]
  wire  _T_25; // @[Misc.scala 209:20]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_30; // @[Misc.scala 213:38]
  wire  _T_31; // @[Misc.scala 213:29]
  wire  _T_34; // @[Misc.scala 209:20]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 212:27]
  wire  _T_45; // @[Misc.scala 213:38]
  wire  _T_46; // @[Misc.scala 213:29]
  wire [3:0] _T_49; // @[Cat.scala 29:58]
  wire [3:0] _T_51; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_300; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_282; // @[OneHot.scala 58:35]
  wire  _T_347; // @[RegisterRouter.scala 59:16]
  wire  _T_349; // @[RegisterRouter.scala 59:16]
  wire  _T_350; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _GEN_24; // @[RegField.scala 134:88]
  wire  _T_154; // @[RegisterRouter.scala 59:16]
  wire  _T_354; // @[RegisterRouter.scala 59:16]
  wire  _T_355; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire  _T_359; // @[RegisterRouter.scala 59:16]
  wire  _T_360; // @[RegisterRouter.scala 59:16]
  wire  _T_207; // @[RegisterRouter.scala 59:16]
  wire  _T_364; // @[RegisterRouter.scala 59:16]
  wire  _T_365; // @[RegisterRouter.scala 59:16]
  wire  _T_230; // @[RegisterRouter.scala 59:16]
  wire  _T_369; // @[RegisterRouter.scala 59:16]
  wire  _T_370; // @[RegisterRouter.scala 59:16]
  wire  _T_253; // @[RegisterRouter.scala 59:16]
  wire  _GEN_62; // @[MuxLiteral.scala 48:10]
  wire  _GEN_63; // @[MuxLiteral.scala 48:10]
  wire  _GEN_64; // @[MuxLiteral.scala 48:10]
  wire  _GEN_65; // @[MuxLiteral.scala 48:10]
  wire  _GEN_66; // @[MuxLiteral.scala 48:10]
  wire  _GEN_67; // @[MuxLiteral.scala 48:10]
  wire  _GEN_77; // @[MuxLiteral.scala 48:10]
  wire  _GEN_68; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_70; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_71; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_72; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_73; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_74; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_75; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_76; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_494; // @[RegisterRouter.scala 59:16]
  wire  _T_495_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_495_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_498; // @[RegisterRouter.scala 65:29]
  LinearSorter lis ( // @[LISDspBlock.scala 55:21]
    .clock(lis_clock),
    .reset(lis_reset),
    .io_in_ready(lis_io_in_ready),
    .io_in_valid(lis_io_in_valid),
    .io_in_bits(lis_io_in_bits),
    .io_lastIn(lis_io_lastIn),
    .io_out_ready(lis_io_out_ready),
    .io_out_valid(lis_io_out_valid),
    .io_out_bits(lis_io_out_bits),
    .io_lastOut(lis_io_lastOut),
    .io_sortedData_0(lis_io_sortedData_0),
    .io_sortedData_1(lis_io_sortedData_1),
    .io_sortedData_2(lis_io_sortedData_2),
    .io_sortedData_3(lis_io_sortedData_3),
    .io_sortedData_4(lis_io_sortedData_4),
    .io_sortedData_5(lis_io_sortedData_5),
    .io_sortedData_6(lis_io_sortedData_6),
    .io_sortedData_7(lis_io_sortedData_7),
    .io_sortedData_8(lis_io_sortedData_8),
    .io_sortedData_9(lis_io_sortedData_9),
    .io_sortedData_10(lis_io_sortedData_10),
    .io_sortedData_11(lis_io_sortedData_11),
    .io_sortedData_12(lis_io_sortedData_12),
    .io_sortedData_13(lis_io_sortedData_13),
    .io_sortedData_14(lis_io_sortedData_14),
    .io_sortedData_15(lis_io_sortedData_15),
    .io_sortedData_16(lis_io_sortedData_16),
    .io_sortedData_17(lis_io_sortedData_17),
    .io_sortedData_18(lis_io_sortedData_18),
    .io_sortedData_19(lis_io_sortedData_19),
    .io_sortedData_20(lis_io_sortedData_20),
    .io_sortedData_21(lis_io_sortedData_21),
    .io_sortedData_22(lis_io_sortedData_22),
    .io_sortedData_23(lis_io_sortedData_23),
    .io_sorterFull(lis_io_sorterFull),
    .io_sorterEmpty(lis_io_sorterEmpty),
    .io_lisSize(lis_io_lisSize)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_stream_in_bits_data; // @[LISDspBlock.scala 71:44]
  assign _GEN_0 = lis_io_sortedData_0; // @[LISDspBlock.scala 92:82]
  assign _GEN_1 = 5'h1 == sendOnOutput ? $signed(lis_io_sortedData_1) : $signed(_GEN_0); // @[LISDspBlock.scala 92:82]
  assign _GEN_2 = 5'h2 == sendOnOutput ? $signed(lis_io_sortedData_2) : $signed(_GEN_1); // @[LISDspBlock.scala 92:82]
  assign _GEN_3 = 5'h3 == sendOnOutput ? $signed(lis_io_sortedData_3) : $signed(_GEN_2); // @[LISDspBlock.scala 92:82]
  assign _GEN_4 = 5'h4 == sendOnOutput ? $signed(lis_io_sortedData_4) : $signed(_GEN_3); // @[LISDspBlock.scala 92:82]
  assign _GEN_5 = 5'h5 == sendOnOutput ? $signed(lis_io_sortedData_5) : $signed(_GEN_4); // @[LISDspBlock.scala 92:82]
  assign _GEN_6 = 5'h6 == sendOnOutput ? $signed(lis_io_sortedData_6) : $signed(_GEN_5); // @[LISDspBlock.scala 92:82]
  assign _GEN_7 = 5'h7 == sendOnOutput ? $signed(lis_io_sortedData_7) : $signed(_GEN_6); // @[LISDspBlock.scala 92:82]
  assign _GEN_8 = 5'h8 == sendOnOutput ? $signed(lis_io_sortedData_8) : $signed(_GEN_7); // @[LISDspBlock.scala 92:82]
  assign _GEN_9 = 5'h9 == sendOnOutput ? $signed(lis_io_sortedData_9) : $signed(_GEN_8); // @[LISDspBlock.scala 92:82]
  assign _GEN_10 = 5'ha == sendOnOutput ? $signed(lis_io_sortedData_10) : $signed(_GEN_9); // @[LISDspBlock.scala 92:82]
  assign _GEN_11 = 5'hb == sendOnOutput ? $signed(lis_io_sortedData_11) : $signed(_GEN_10); // @[LISDspBlock.scala 92:82]
  assign _GEN_12 = 5'hc == sendOnOutput ? $signed(lis_io_sortedData_12) : $signed(_GEN_11); // @[LISDspBlock.scala 92:82]
  assign _GEN_13 = 5'hd == sendOnOutput ? $signed(lis_io_sortedData_13) : $signed(_GEN_12); // @[LISDspBlock.scala 92:82]
  assign _GEN_14 = 5'he == sendOnOutput ? $signed(lis_io_sortedData_14) : $signed(_GEN_13); // @[LISDspBlock.scala 92:82]
  assign _GEN_15 = 5'hf == sendOnOutput ? $signed(lis_io_sortedData_15) : $signed(_GEN_14); // @[LISDspBlock.scala 92:82]
  assign _GEN_16 = 5'h10 == sendOnOutput ? $signed(lis_io_sortedData_16) : $signed(_GEN_15); // @[LISDspBlock.scala 92:82]
  assign _GEN_17 = 5'h11 == sendOnOutput ? $signed(lis_io_sortedData_17) : $signed(_GEN_16); // @[LISDspBlock.scala 92:82]
  assign _GEN_18 = 5'h12 == sendOnOutput ? $signed(lis_io_sortedData_18) : $signed(_GEN_17); // @[LISDspBlock.scala 92:82]
  assign _GEN_19 = 5'h13 == sendOnOutput ? $signed(lis_io_sortedData_19) : $signed(_GEN_18); // @[LISDspBlock.scala 92:82]
  assign _GEN_20 = 5'h14 == sendOnOutput ? $signed(lis_io_sortedData_20) : $signed(_GEN_19); // @[LISDspBlock.scala 92:82]
  assign _GEN_21 = 5'h15 == sendOnOutput ? $signed(lis_io_sortedData_21) : $signed(_GEN_20); // @[LISDspBlock.scala 92:82]
  assign _GEN_22 = 5'h16 == sendOnOutput ? $signed(lis_io_sortedData_22) : $signed(_GEN_21); // @[LISDspBlock.scala 92:82]
  assign _T_4 = 5'h17 == sendOnOutput ? $signed(lis_io_sortedData_23) : $signed(_GEN_22); // @[LISDspBlock.scala 92:82]
  assign _T_7 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_8 = auto_mem_in_ar_valid | _T_7; // @[RegisterRouter.scala 40:26]
  assign _T_9 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_52_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_16 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_281 = {_T_16[4],_T_16[3],_T_16[2]}; // @[Cat.scala 29:58]
  assign _T_56 = _T_16[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_64 = _T_56 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_10 = _T_52_ready & _T_9; // @[RegisterRouter.scala 42:26]
  assign _T_19 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_21 = _T_19 | 2'h1; // @[Misc.scala 200:81]
  assign _T_22 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_25 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_27 = _T_21[1] & _T_25; // @[Misc.scala 213:38]
  assign _T_28 = _T_22 | _T_27; // @[Misc.scala 213:29]
  assign _T_30 = _T_21[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_31 = _T_22 | _T_30; // @[Misc.scala 213:29]
  assign _T_34 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_35 = _T_25 & _T_34; // @[Misc.scala 212:27]
  assign _T_36 = _T_21[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = _T_25 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_39 = _T_21[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & _T_34; // @[Misc.scala 212:27]
  assign _T_42 = _T_21[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_31 | _T_42; // @[Misc.scala 213:29]
  assign _T_44 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_45 = _T_21[0] & _T_44; // @[Misc.scala 213:38]
  assign _T_46 = _T_31 | _T_45; // @[Misc.scala 213:29]
  assign _T_49 = {_T_46,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  assign _T_51 = auto_mem_in_ar_valid ? _T_49 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_51[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_51[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_51[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_51[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_300 = _T_8 & _T_52_ready; // @[RegisterRouter.scala 59:16]
  assign _T_282 = 8'h1 << _T_281; // @[OneHot.scala 58:35]
  assign _T_347 = _T_300 & _T_9; // @[RegisterRouter.scala 59:16]
  assign _T_349 = _T_347 & _T_282[0]; // @[RegisterRouter.scala 59:16]
  assign _T_350 = _T_349 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_350 & _T_89[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_24 = _T_115 ? auto_mem_in_w_bits_data[0] : sortDir; // @[RegField.scala 134:88]
  assign _T_154 = _T_89[4:0] == 5'h1f; // @[RegisterRouter.scala 59:16]
  assign _T_354 = _T_347 & _T_282[1]; // @[RegisterRouter.scala 59:16]
  assign _T_355 = _T_354 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_355 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _T_359 = _T_347 & _T_282[2]; // @[RegisterRouter.scala 59:16]
  assign _T_360 = _T_359 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_207 = _T_360 & _T_89[0]; // @[RegisterRouter.scala 59:16]
  assign _T_364 = _T_347 & _T_282[3]; // @[RegisterRouter.scala 59:16]
  assign _T_365 = _T_364 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_230 = _T_365 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _T_369 = _T_347 & _T_282[4]; // @[RegisterRouter.scala 59:16]
  assign _T_370 = _T_369 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_253 = _T_370 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _GEN_62 = 3'h1 == _T_281 ? _T_64 : _T_64; // @[MuxLiteral.scala 48:10]
  assign _GEN_63 = 3'h2 == _T_281 ? _T_64 : _GEN_62; // @[MuxLiteral.scala 48:10]
  assign _GEN_64 = 3'h3 == _T_281 ? _T_64 : _GEN_63; // @[MuxLiteral.scala 48:10]
  assign _GEN_65 = 3'h4 == _T_281 ? _T_64 : _GEN_64; // @[MuxLiteral.scala 48:10]
  assign _GEN_66 = 3'h5 == _T_281 ? _T_64 : _GEN_65; // @[MuxLiteral.scala 48:10]
  assign _GEN_67 = 3'h6 == _T_281 ? _T_64 : _GEN_66; // @[MuxLiteral.scala 48:10]
  assign _GEN_77 = 3'h7 == _T_281; // @[MuxLiteral.scala 48:10]
  assign _GEN_68 = _GEN_77 | _GEN_67; // @[MuxLiteral.scala 48:10]
  assign _T_492_0 = {{4'd0}, sortDir}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_70 = 3'h1 == _T_281 ? lisSize : _T_492_0; // @[MuxLiteral.scala 48:10]
  assign _T_492_2 = {{4'd0}, flushData}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_71 = 3'h2 == _T_281 ? _T_492_2 : _GEN_70; // @[MuxLiteral.scala 48:10]
  assign _GEN_72 = 3'h3 == _T_281 ? discardPos : _GEN_71; // @[MuxLiteral.scala 48:10]
  assign _GEN_73 = 3'h4 == _T_281 ? sendOnOutput : _GEN_72; // @[MuxLiteral.scala 48:10]
  assign _T_492_5 = {{4'd0}, sorterFull}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_74 = 3'h5 == _T_281 ? _T_492_5 : _GEN_73; // @[MuxLiteral.scala 48:10]
  assign _T_492_6 = {{4'd0}, sorterEmpty}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_75 = 3'h6 == _T_281 ? _T_492_6 : _GEN_74; // @[MuxLiteral.scala 48:10]
  assign _GEN_76 = 3'h7 == _T_281 ? 5'h0 : _GEN_75; // @[MuxLiteral.scala 48:10]
  assign _T_494 = _GEN_68 ? _GEN_76 : 5'h0; // @[RegisterRouter.scala 59:16]
  assign _T_495_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_495_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_498 = ~_T_495_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_10 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_10 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_495_valid & _T_498; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_495_valid & _T_495_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = lis_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = lis_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {lis_io_out_bits,_T_4}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = lis_io_lastOut; // @[LazyModule.scala 173:49]
  assign lis_clock = clock;
  assign lis_reset = reset;
  assign lis_io_in_valid = auto_stream_in_valid; // @[LISDspBlock.scala 70:21]
  assign lis_io_in_bits = _T_2[15:0]; // @[LISDspBlock.scala 71:20]
  assign lis_io_lastIn = auto_stream_in_bits_last; // @[LISDspBlock.scala 69:19]
  assign lis_io_out_ready = auto_stream_out_ready; // @[LISDspBlock.scala 91:22]
  assign lis_io_lisSize = {{1'd0}, lisSize}; // @[LISDspBlock.scala 79:26]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_7; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{27'd0}, _T_494}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_495_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sortDir = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flushData = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  discardPos = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sendOnOutput = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  lisSize = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sorterFull = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sorterEmpty = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sortDir <= reset | _GEN_24;
    if (reset) begin
      flushData <= 1'h0;
    end else if (_T_207) begin
      flushData <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      discardPos <= 5'h0;
    end else if (_T_230) begin
      discardPos <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      sendOnOutput <= 5'h0;
    end else if (_T_253) begin
      sendOnOutput <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      lisSize <= 5'h18;
    end else if (_T_161) begin
      lisSize <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      sorterFull <= 1'h0;
    end else begin
      sorterFull <= lis_io_sorterFull;
    end
    sorterEmpty <= reset | lis_io_sorterEmpty;
  end
endmodule
module AXI4StreamMux(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_4_ready,
  input         auto_stream_in_4_valid,
  input  [31:0] auto_stream_in_4_bits_data,
  input         auto_stream_in_4_bits_last,
  output        auto_stream_in_3_ready,
  input         auto_stream_in_3_valid,
  input  [31:0] auto_stream_in_3_bits_data,
  input         auto_stream_in_3_bits_last,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _GEN_35; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _GEN_44; // @[Mux.scala 45:41]
  wire  _T_8; // @[Mux.scala 40:46]
  wire [2:0] _T_10; // @[Mux.scala 41:29]
  wire  _T_11; // @[Mux.scala 45:28]
  wire  _T_12; // @[Mux.scala 45:28]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _T_14; // @[Mux.scala 45:28]
  wire  _T_15; // @[Mux.scala 45:28]
  wire  _T_17; // @[RegisterRouter.scala 40:39]
  wire  _T_18; // @[RegisterRouter.scala 40:26]
  wire  _T_19; // @[RegisterRouter.scala 42:29]
  wire  _T_62_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_26; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_66; // @[RegisterRouter.scala 59:16]
  wire  _T_68; // @[RegisterRouter.scala 59:16]
  wire  _T_20; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_29; // @[OneHot.scala 65:12]
  wire [1:0] _T_31; // @[Misc.scala 200:81]
  wire  _T_32; // @[Misc.scala 204:21]
  wire  _T_35; // @[Misc.scala 209:20]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 213:38]
  wire  _T_41; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 209:20]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire  _T_54; // @[Misc.scala 212:27]
  wire  _T_55; // @[Misc.scala 213:38]
  wire  _T_56; // @[Misc.scala 213:29]
  wire [3:0] _T_59; // @[Cat.scala 29:58]
  wire [3:0] _T_61; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_108; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_155; // @[OneHot.scala 58:35]
  wire  _T_178; // @[RegisterRouter.scala 59:16]
  wire  _T_185; // @[RegisterRouter.scala 59:16]
  wire  _T_186; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_180; // @[RegisterRouter.scala 59:16]
  wire  _T_181; // @[RegisterRouter.scala 59:16]
  wire  _T_138; // @[RegisterRouter.scala 59:16]
  wire  _GEN_101; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_103; // @[MuxLiteral.scala 48:10]
  wire [2:0] _T_235; // @[RegisterRouter.scala 59:16]
  wire  _T_236_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_236_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_239; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? auto_stream_in_3_bits_last : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? auto_stream_in_3_bits_data : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 ? auto_stream_in_3_valid : _GEN_25; // @[Mux.scala 45:41]
  assign _GEN_35 = _T_6 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _GEN_44 = _T_7 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_8 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_10 = _T_8 ? 3'h5 : sels_1; // @[Mux.scala 41:29]
  assign _T_11 = _T_10 == 3'h0; // @[Mux.scala 45:28]
  assign _T_12 = _T_10 == 3'h1; // @[Mux.scala 45:28]
  assign _T_13 = _T_10 == 3'h2; // @[Mux.scala 45:28]
  assign _T_14 = _T_10 == 3'h3; // @[Mux.scala 45:28]
  assign _T_15 = _T_10 == 3'h4; // @[Mux.scala 45:28]
  assign _T_17 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_18 = auto_register_in_ar_valid | _T_17; // @[RegisterRouter.scala 40:26]
  assign _T_19 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_62_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_26 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_66 = _T_26[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_68 = _T_66 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_20 = _T_62_ready & _T_19; // @[RegisterRouter.scala 42:26]
  assign _T_29 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_31 = _T_29 | 2'h1; // @[Misc.scala 200:81]
  assign _T_32 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_35 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_37 = _T_31[1] & _T_35; // @[Misc.scala 213:38]
  assign _T_38 = _T_32 | _T_37; // @[Misc.scala 213:29]
  assign _T_40 = _T_31[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_41 = _T_32 | _T_40; // @[Misc.scala 213:29]
  assign _T_44 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_45 = _T_35 & _T_44; // @[Misc.scala 212:27]
  assign _T_46 = _T_31[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_38 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = _T_35 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_49 = _T_31[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_register_in_ar_bits_addr[1] & _T_44; // @[Misc.scala 212:27]
  assign _T_52 = _T_31[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_41 | _T_52; // @[Misc.scala 213:29]
  assign _T_54 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_55 = _T_31[0] & _T_54; // @[Misc.scala 213:38]
  assign _T_56 = _T_41 | _T_55; // @[Misc.scala 213:29]
  assign _T_59 = {_T_56,_T_53,_T_50,_T_47}; // @[Cat.scala 29:58]
  assign _T_61 = auto_register_in_ar_valid ? _T_59 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_61[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_61[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_61[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_61[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_108 = _T_89[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_18 & _T_62_ready; // @[RegisterRouter.scala 59:16]
  assign _T_155 = 2'h1 << _T_26[2]; // @[OneHot.scala 58:35]
  assign _T_178 = _T_161 & _T_19; // @[RegisterRouter.scala 59:16]
  assign _T_185 = _T_178 & _T_155[1]; // @[RegisterRouter.scala 59:16]
  assign _T_186 = _T_185 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_186 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _T_180 = _T_178 & _T_155[0]; // @[RegisterRouter.scala 59:16]
  assign _T_181 = _T_180 & _T_68; // @[RegisterRouter.scala 59:16]
  assign _T_138 = _T_181 & _T_108; // @[RegisterRouter.scala 59:16]
  assign _GEN_101 = _T_26[2] ? _T_68 : _T_68; // @[MuxLiteral.scala 48:10]
  assign _GEN_103 = _T_26[2] ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _T_235 = _GEN_101 ? _GEN_103 : 3'h0; // @[RegisterRouter.scala 59:16]
  assign _T_236_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_236_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_239 = ~_T_236_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_20 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_20 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_236_valid & _T_239; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_236_valid & _T_236_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_4_ready = _T_15 | _GEN_44; // @[LazyModule.scala 173:31]
  assign auto_stream_in_3_ready = _T_14 | _GEN_35; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_13 | _GEN_26; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_12 | _GEN_17; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_11 | _GEN_8; // @[LazyModule.scala 173:31]
  assign auto_stream_out_0_valid = _T_7 ? auto_stream_in_4_valid : _GEN_34; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_7 ? auto_stream_in_4_bits_data : _GEN_33; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_7 ? auto_stream_in_4_bits_last : _GEN_30; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_17; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _T_235}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_236_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h5;
    end else if (_T_138) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h5;
    end else if (_T_115) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module PE_24(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_rightOutData,
  output        io_currDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_rightOutData = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = 1'h1; // @[PE.scala 56:30]
  assign ctrlLogic_io_rightCompOut = _T_3 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_3 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= 16'sh0;
      end else begin
        saveCellData <= io_rightNBR_data;
      end
    end
  end
endmodule
module PE_25(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_26(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_27(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_28(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_29(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_30(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_31(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_32(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_33(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_34(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_35(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_36(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_37(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_38(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_39(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_40(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_41(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_42(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_43(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_44(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_45(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_46(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  input  [15:0] io_rightNBR_data,
  input         io_rightNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  input         io_rightPropDiscard,
  output [15:0] io_leftOutData,
  output [15:0] io_rightOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  _T_3; // @[PE.scala 62:40]
  wire  _T_4; // @[PE.scala 62:37]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  wire [15:0] _T_20; // @[PE.scala 147:27]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign _T_3 = ~io_lastCell; // @[PE.scala 62:40]
  assign _T_4 = io_active & _T_3; // @[PE.scala 62:37]
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign _T_20 = compRes ? $signed(io_inData) : $signed(saveCellData); // @[PE.scala 147:27]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_rightOutData = io_active ? $signed(_T_20) : $signed(saveCellData); // @[PE.scala 147:21 PE.scala 150:21]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = _T_4 & io_rightNBR_compRes; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = _T_4 & io_rightPropDiscard; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= io_rightNBR_data;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module PE_47(
  input         clock,
  input         reset,
  input         io_enableSort,
  input  [1:0]  io_state,
  input  [15:0] io_leftNBR_data,
  input         io_leftNBR_compRes,
  output [15:0] io_currCell_data,
  output        io_currCell_compRes,
  input         io_lastCell,
  input         io_active,
  input         io_discard,
  input  [15:0] io_inData,
  output [15:0] io_leftOutData,
  output        io_currDiscard,
  output        io_toLeftPropDiscard
);
  wire  ctrlLogic_io_currCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightCompOut; // @[PE.scala 53:25]
  wire  ctrlLogic_io_currDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rightPropDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_propDiscard; // @[PE.scala 53:25]
  wire  ctrlLogic_io_load; // @[PE.scala 53:25]
  wire  ctrlLogic_io_leftRightShift; // @[PE.scala 53:25]
  wire  ctrlLogic_io_rstPEregs; // @[PE.scala 53:25]
  wire  load; // @[PE.scala 89:29]
  reg [15:0] saveCellData; // @[PE.scala 112:29]
  reg [31:0] _RAND_0;
  wire  _T_9; // @[PE.scala 114:18]
  wire  compRes; // @[FixedPointTypeClass.scala 53:59]
  PEControlLogic ctrlLogic ( // @[PE.scala 53:25]
    .io_currCompOut(ctrlLogic_io_currCompOut),
    .io_leftCompOut(ctrlLogic_io_leftCompOut),
    .io_rightCompOut(ctrlLogic_io_rightCompOut),
    .io_currDiscard(ctrlLogic_io_currDiscard),
    .io_rightPropDiscard(ctrlLogic_io_rightPropDiscard),
    .io_propDiscard(ctrlLogic_io_propDiscard),
    .io_load(ctrlLogic_io_load),
    .io_leftRightShift(ctrlLogic_io_leftRightShift),
    .io_rstPEregs(ctrlLogic_io_rstPEregs)
  );
  assign load = io_enableSort & ctrlLogic_io_load; // @[PE.scala 89:29]
  assign _T_9 = io_state == 2'h0; // @[PE.scala 114:18]
  assign compRes = $signed(saveCellData) < $signed(io_inData); // @[FixedPointTypeClass.scala 53:59]
  assign io_currCell_data = saveCellData; // @[PE.scala 137:20]
  assign io_currCell_compRes = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 136:23]
  assign io_leftOutData = compRes ? $signed(saveCellData) : $signed(io_inData); // @[PE.scala 143:20]
  assign io_currDiscard = io_discard; // @[PE.scala 168:20]
  assign io_toLeftPropDiscard = ctrlLogic_io_propDiscard; // @[PE.scala 133:26]
  assign ctrlLogic_io_currCompOut = $signed(saveCellData) < $signed(io_inData); // @[PE.scala 126:28]
  assign ctrlLogic_io_leftCompOut = io_leftNBR_compRes; // @[PE.scala 59:30]
  assign ctrlLogic_io_rightCompOut = 1'h0; // @[PE.scala 63:31 PE.scala 67:31]
  assign ctrlLogic_io_currDiscard = io_discard; // @[PE.scala 167:30]
  assign ctrlLogic_io_rightPropDiscard = 1'h0; // @[PE.scala 64:35 PE.scala 68:35]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saveCellData = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      saveCellData <= -16'sh8000;
    end else if (_T_9) begin
      saveCellData <= -16'sh8000;
    end else if (load) begin
      if (io_lastCell) begin
        saveCellData <= io_leftNBR_data;
      end else if (io_active) begin
        if (ctrlLogic_io_leftRightShift) begin
          saveCellData <= 16'sh0;
        end else begin
          saveCellData <= io_leftNBR_data;
        end
      end else begin
        saveCellData <= -16'sh8000;
      end
    end
  end
endmodule
module LinearSorter_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut,
  output [15:0] io_sortedData_0,
  output [15:0] io_sortedData_1,
  output [15:0] io_sortedData_2,
  output [15:0] io_sortedData_3,
  output [15:0] io_sortedData_4,
  output [15:0] io_sortedData_5,
  output [15:0] io_sortedData_6,
  output [15:0] io_sortedData_7,
  output [15:0] io_sortedData_8,
  output [15:0] io_sortedData_9,
  output [15:0] io_sortedData_10,
  output [15:0] io_sortedData_11,
  output [15:0] io_sortedData_12,
  output [15:0] io_sortedData_13,
  output [15:0] io_sortedData_14,
  output [15:0] io_sortedData_15,
  output [15:0] io_sortedData_16,
  output [15:0] io_sortedData_17,
  output [15:0] io_sortedData_18,
  output [15:0] io_sortedData_19,
  output [15:0] io_sortedData_20,
  output [15:0] io_sortedData_21,
  output [15:0] io_sortedData_22,
  output [15:0] io_sortedData_23,
  output        io_sorterFull,
  output        io_sorterEmpty,
  input  [5:0]  io_lisSize,
  input  [4:0]  io_discardPos
);
  wire  PEChain_0_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_0_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_1_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_2_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_3_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_4_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_5_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_6_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_7_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_8_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_9_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_10_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_11_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_12_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_13_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_14_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_15_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_16_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_17_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_18_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_19_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_20_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_21_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_22_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_23_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_inData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  reg  initialInDone; // @[LinearSorter.scala 67:30]
  reg [31:0] _RAND_0;
  reg [4:0] cntInData; // @[LinearSorter.scala 68:26]
  reg [31:0] _RAND_1;
  reg [1:0] state; // @[LinearSorter.scala 78:22]
  reg [31:0] _RAND_2;
  reg [5:0] lisSizeReg; // @[LinearSorter.scala 81:27]
  reg [31:0] _RAND_3;
  wire [5:0] _T_1; // @[LinearSorter.scala 86:43]
  wire  _T_96; // @[Decoupled.scala 40:37]
  wire [4:0] _T_98; // @[LinearSorter.scala 92:28]
  wire  _T_99; // @[LinearSorter.scala 94:20]
  wire [5:0] _GEN_111; // @[LinearSorter.scala 98:19]
  wire  _T_102; // @[LinearSorter.scala 98:19]
  wire  _T_104; // @[LinearSorter.scala 98:42]
  wire  _T_113; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_7; // @[LinearSorter.scala 117:27]
  wire  _T_115; // @[Conditional.scala 37:30]
  wire  fireLastIn; // @[LinearSorter.scala 111:30]
  wire [1:0] _GEN_8; // @[LinearSorter.scala 120:62]
  wire  _T_117; // @[Conditional.scala 37:30]
  reg [4:0] cntOutData; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_4;
  wire [5:0] _GEN_112; // @[LinearSorter.scala 125:28]
  wire  _T_120; // @[LinearSorter.scala 125:28]
  wire [1:0] _GEN_9; // @[LinearSorter.scala 125:50]
  wire [1:0] _GEN_10; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_11; // @[Conditional.scala 39:67]
  wire [1:0] state_next; // @[Conditional.scala 40:58]
  wire  _T_105; // @[LinearSorter.scala 101:25]
  wire  _GEN_2; // @[LinearSorter.scala 101:36]
  wire  _GEN_3; // @[LinearSorter.scala 98:59]
  wire  _T_106; // @[LinearSorter.scala 106:29]
  wire  _T_107; // @[LinearSorter.scala 106:54]
  wire  enable; // @[LinearSorter.scala 106:45]
  wire  _T_109; // @[LISutil.scala 13:24]
  wire [4:0] _T_111; // @[LISutil.scala 14:22]
  wire  _T_121; // @[LinearSorter.scala 137:33]
  wire [15:0] outputData_0; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] outputData_1; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_16; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_2; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_17; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_3; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_18; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_4; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_19; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_5; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_20; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_6; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_21; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_7; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_22; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_8; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_23; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_9; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_24; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_10; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_25; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_11; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_26; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_12; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_27; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_13; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_28; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_14; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_29; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_15; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_30; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_16; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_31; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_17; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_32; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_18; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_33; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_19; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_34; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_20; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_35; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_21; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_36; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_22; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_37; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_23; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_38; // @[LinearSorter.scala 137:21]
  wire  _T_132; // @[LinearSorter.scala 160:26]
  wire  _GEN_39; // @[LinearSorter.scala 160:80]
  wire  _T_136; // @[LinearSorter.scala 168:63]
  wire  _T_142; // @[LinearSorter.scala 160:26]
  wire  _GEN_41; // @[LinearSorter.scala 160:80]
  wire  _T_152; // @[LinearSorter.scala 160:26]
  wire  _GEN_43; // @[LinearSorter.scala 160:80]
  wire  _T_162; // @[LinearSorter.scala 160:26]
  wire  _GEN_45; // @[LinearSorter.scala 160:80]
  wire  _T_172; // @[LinearSorter.scala 160:26]
  wire  _GEN_47; // @[LinearSorter.scala 160:80]
  wire  _T_182; // @[LinearSorter.scala 160:26]
  wire  _GEN_49; // @[LinearSorter.scala 160:80]
  wire  _T_192; // @[LinearSorter.scala 160:26]
  wire  _GEN_51; // @[LinearSorter.scala 160:80]
  wire  _T_202; // @[LinearSorter.scala 160:26]
  wire  _GEN_53; // @[LinearSorter.scala 160:80]
  wire  _T_212; // @[LinearSorter.scala 160:26]
  wire  _GEN_55; // @[LinearSorter.scala 160:80]
  wire  _T_222; // @[LinearSorter.scala 160:26]
  wire  _GEN_57; // @[LinearSorter.scala 160:80]
  wire  _T_232; // @[LinearSorter.scala 160:26]
  wire  _GEN_59; // @[LinearSorter.scala 160:80]
  wire  _T_242; // @[LinearSorter.scala 160:26]
  wire  _GEN_61; // @[LinearSorter.scala 160:80]
  wire  _T_252; // @[LinearSorter.scala 160:26]
  wire  _GEN_63; // @[LinearSorter.scala 160:80]
  wire  _T_262; // @[LinearSorter.scala 160:26]
  wire  _GEN_65; // @[LinearSorter.scala 160:80]
  wire  _T_272; // @[LinearSorter.scala 160:26]
  wire  _GEN_67; // @[LinearSorter.scala 160:80]
  wire  _T_282; // @[LinearSorter.scala 160:26]
  wire  _GEN_69; // @[LinearSorter.scala 160:80]
  wire  _T_292; // @[LinearSorter.scala 160:26]
  wire  _GEN_71; // @[LinearSorter.scala 160:80]
  wire  _T_302; // @[LinearSorter.scala 160:26]
  wire  _GEN_73; // @[LinearSorter.scala 160:80]
  wire  _T_312; // @[LinearSorter.scala 160:26]
  wire  _GEN_75; // @[LinearSorter.scala 160:80]
  wire  _T_322; // @[LinearSorter.scala 160:26]
  wire  _GEN_77; // @[LinearSorter.scala 160:80]
  wire  _T_332; // @[LinearSorter.scala 160:26]
  wire  _GEN_79; // @[LinearSorter.scala 160:80]
  wire  _T_342; // @[LinearSorter.scala 160:26]
  wire  _GEN_81; // @[LinearSorter.scala 160:80]
  wire  _T_352; // @[LinearSorter.scala 160:26]
  wire  _GEN_83; // @[LinearSorter.scala 160:80]
  wire  _T_362; // @[LinearSorter.scala 160:26]
  wire  _GEN_85; // @[LinearSorter.scala 160:80]
  wire  discardSignals_2; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_1; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_0; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_5; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_4; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_3; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [5:0] _T_372; // @[LinearSorter.scala 177:50]
  wire  discardSignals_8; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_7; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_6; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_11; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_10; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_9; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [11:0] _T_378; // @[LinearSorter.scala 177:50]
  wire  discardSignals_14; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_13; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_12; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_17; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_16; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_15; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [5:0] _T_383; // @[LinearSorter.scala 177:50]
  wire  discardSignals_20; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_19; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_18; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_23; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_22; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_21; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [23:0] _T_390; // @[LinearSorter.scala 177:50]
  wire [4:0] _T_415; // @[Mux.scala 47:69]
  wire [4:0] _T_416; // @[Mux.scala 47:69]
  wire [4:0] _T_417; // @[Mux.scala 47:69]
  wire [4:0] _T_418; // @[Mux.scala 47:69]
  wire [4:0] _T_419; // @[Mux.scala 47:69]
  wire [4:0] _T_420; // @[Mux.scala 47:69]
  wire [4:0] _T_421; // @[Mux.scala 47:69]
  wire [4:0] _T_422; // @[Mux.scala 47:69]
  wire [4:0] _T_423; // @[Mux.scala 47:69]
  wire [4:0] _T_424; // @[Mux.scala 47:69]
  wire [4:0] _T_425; // @[Mux.scala 47:69]
  wire [4:0] _T_426; // @[Mux.scala 47:69]
  wire [4:0] _T_427; // @[Mux.scala 47:69]
  wire [4:0] _T_428; // @[Mux.scala 47:69]
  wire [4:0] _T_429; // @[Mux.scala 47:69]
  wire [4:0] _T_430; // @[Mux.scala 47:69]
  wire [4:0] _T_431; // @[Mux.scala 47:69]
  wire [4:0] _T_432; // @[Mux.scala 47:69]
  wire [4:0] _T_433; // @[Mux.scala 47:69]
  wire [4:0] _T_434; // @[Mux.scala 47:69]
  wire [4:0] _T_435; // @[Mux.scala 47:69]
  wire [4:0] _T_436; // @[Mux.scala 47:69]
  wire [4:0] getDiscarded; // @[Mux.scala 47:69]
  wire  _T_438; // @[LinearSorter.scala 199:49]
  wire [15:0] _GEN_88; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_89; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_90; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_91; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_92; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_93; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_94; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_95; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_96; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_97; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_98; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_99; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_100; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_101; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_102; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_103; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_104; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_105; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_106; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_107; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_108; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_109; // @[LinearSorter.scala 206:15]
  wire  _T_444; // @[LinearSorter.scala 208:18]
  wire  _T_446; // @[LinearSorter.scala 208:49]
  wire  _T_448; // @[LinearSorter.scala 209:33]
  PE_24 PEChain_0 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_0_clock),
    .reset(PEChain_0_reset),
    .io_enableSort(PEChain_0_io_enableSort),
    .io_state(PEChain_0_io_state),
    .io_rightNBR_data(PEChain_0_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_0_io_rightNBR_compRes),
    .io_currCell_data(PEChain_0_io_currCell_data),
    .io_currCell_compRes(PEChain_0_io_currCell_compRes),
    .io_lastCell(PEChain_0_io_lastCell),
    .io_discard(PEChain_0_io_discard),
    .io_inData(PEChain_0_io_inData),
    .io_rightPropDiscard(PEChain_0_io_rightPropDiscard),
    .io_rightOutData(PEChain_0_io_rightOutData),
    .io_currDiscard(PEChain_0_io_currDiscard)
  );
  PE_25 PEChain_1 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_1_clock),
    .reset(PEChain_1_reset),
    .io_enableSort(PEChain_1_io_enableSort),
    .io_state(PEChain_1_io_state),
    .io_leftNBR_data(PEChain_1_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_1_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_1_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_1_io_rightNBR_compRes),
    .io_currCell_data(PEChain_1_io_currCell_data),
    .io_currCell_compRes(PEChain_1_io_currCell_compRes),
    .io_lastCell(PEChain_1_io_lastCell),
    .io_active(PEChain_1_io_active),
    .io_discard(PEChain_1_io_discard),
    .io_inData(PEChain_1_io_inData),
    .io_rightPropDiscard(PEChain_1_io_rightPropDiscard),
    .io_leftOutData(PEChain_1_io_leftOutData),
    .io_rightOutData(PEChain_1_io_rightOutData),
    .io_currDiscard(PEChain_1_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_1_io_toLeftPropDiscard)
  );
  PE_26 PEChain_2 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_2_clock),
    .reset(PEChain_2_reset),
    .io_enableSort(PEChain_2_io_enableSort),
    .io_state(PEChain_2_io_state),
    .io_leftNBR_data(PEChain_2_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_2_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_2_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_2_io_rightNBR_compRes),
    .io_currCell_data(PEChain_2_io_currCell_data),
    .io_currCell_compRes(PEChain_2_io_currCell_compRes),
    .io_lastCell(PEChain_2_io_lastCell),
    .io_active(PEChain_2_io_active),
    .io_discard(PEChain_2_io_discard),
    .io_inData(PEChain_2_io_inData),
    .io_rightPropDiscard(PEChain_2_io_rightPropDiscard),
    .io_leftOutData(PEChain_2_io_leftOutData),
    .io_rightOutData(PEChain_2_io_rightOutData),
    .io_currDiscard(PEChain_2_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_2_io_toLeftPropDiscard)
  );
  PE_27 PEChain_3 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_3_clock),
    .reset(PEChain_3_reset),
    .io_enableSort(PEChain_3_io_enableSort),
    .io_state(PEChain_3_io_state),
    .io_leftNBR_data(PEChain_3_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_3_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_3_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_3_io_rightNBR_compRes),
    .io_currCell_data(PEChain_3_io_currCell_data),
    .io_currCell_compRes(PEChain_3_io_currCell_compRes),
    .io_lastCell(PEChain_3_io_lastCell),
    .io_active(PEChain_3_io_active),
    .io_discard(PEChain_3_io_discard),
    .io_inData(PEChain_3_io_inData),
    .io_rightPropDiscard(PEChain_3_io_rightPropDiscard),
    .io_leftOutData(PEChain_3_io_leftOutData),
    .io_rightOutData(PEChain_3_io_rightOutData),
    .io_currDiscard(PEChain_3_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_3_io_toLeftPropDiscard)
  );
  PE_28 PEChain_4 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_4_clock),
    .reset(PEChain_4_reset),
    .io_enableSort(PEChain_4_io_enableSort),
    .io_state(PEChain_4_io_state),
    .io_leftNBR_data(PEChain_4_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_4_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_4_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_4_io_rightNBR_compRes),
    .io_currCell_data(PEChain_4_io_currCell_data),
    .io_currCell_compRes(PEChain_4_io_currCell_compRes),
    .io_lastCell(PEChain_4_io_lastCell),
    .io_active(PEChain_4_io_active),
    .io_discard(PEChain_4_io_discard),
    .io_inData(PEChain_4_io_inData),
    .io_rightPropDiscard(PEChain_4_io_rightPropDiscard),
    .io_leftOutData(PEChain_4_io_leftOutData),
    .io_rightOutData(PEChain_4_io_rightOutData),
    .io_currDiscard(PEChain_4_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_4_io_toLeftPropDiscard)
  );
  PE_29 PEChain_5 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_5_clock),
    .reset(PEChain_5_reset),
    .io_enableSort(PEChain_5_io_enableSort),
    .io_state(PEChain_5_io_state),
    .io_leftNBR_data(PEChain_5_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_5_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_5_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_5_io_rightNBR_compRes),
    .io_currCell_data(PEChain_5_io_currCell_data),
    .io_currCell_compRes(PEChain_5_io_currCell_compRes),
    .io_lastCell(PEChain_5_io_lastCell),
    .io_active(PEChain_5_io_active),
    .io_discard(PEChain_5_io_discard),
    .io_inData(PEChain_5_io_inData),
    .io_rightPropDiscard(PEChain_5_io_rightPropDiscard),
    .io_leftOutData(PEChain_5_io_leftOutData),
    .io_rightOutData(PEChain_5_io_rightOutData),
    .io_currDiscard(PEChain_5_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_5_io_toLeftPropDiscard)
  );
  PE_30 PEChain_6 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_6_clock),
    .reset(PEChain_6_reset),
    .io_enableSort(PEChain_6_io_enableSort),
    .io_state(PEChain_6_io_state),
    .io_leftNBR_data(PEChain_6_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_6_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_6_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_6_io_rightNBR_compRes),
    .io_currCell_data(PEChain_6_io_currCell_data),
    .io_currCell_compRes(PEChain_6_io_currCell_compRes),
    .io_lastCell(PEChain_6_io_lastCell),
    .io_active(PEChain_6_io_active),
    .io_discard(PEChain_6_io_discard),
    .io_inData(PEChain_6_io_inData),
    .io_rightPropDiscard(PEChain_6_io_rightPropDiscard),
    .io_leftOutData(PEChain_6_io_leftOutData),
    .io_rightOutData(PEChain_6_io_rightOutData),
    .io_currDiscard(PEChain_6_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_6_io_toLeftPropDiscard)
  );
  PE_31 PEChain_7 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_7_clock),
    .reset(PEChain_7_reset),
    .io_enableSort(PEChain_7_io_enableSort),
    .io_state(PEChain_7_io_state),
    .io_leftNBR_data(PEChain_7_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_7_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_7_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_7_io_rightNBR_compRes),
    .io_currCell_data(PEChain_7_io_currCell_data),
    .io_currCell_compRes(PEChain_7_io_currCell_compRes),
    .io_lastCell(PEChain_7_io_lastCell),
    .io_active(PEChain_7_io_active),
    .io_discard(PEChain_7_io_discard),
    .io_inData(PEChain_7_io_inData),
    .io_rightPropDiscard(PEChain_7_io_rightPropDiscard),
    .io_leftOutData(PEChain_7_io_leftOutData),
    .io_rightOutData(PEChain_7_io_rightOutData),
    .io_currDiscard(PEChain_7_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_7_io_toLeftPropDiscard)
  );
  PE_32 PEChain_8 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_8_clock),
    .reset(PEChain_8_reset),
    .io_enableSort(PEChain_8_io_enableSort),
    .io_state(PEChain_8_io_state),
    .io_leftNBR_data(PEChain_8_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_8_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_8_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_8_io_rightNBR_compRes),
    .io_currCell_data(PEChain_8_io_currCell_data),
    .io_currCell_compRes(PEChain_8_io_currCell_compRes),
    .io_lastCell(PEChain_8_io_lastCell),
    .io_active(PEChain_8_io_active),
    .io_discard(PEChain_8_io_discard),
    .io_inData(PEChain_8_io_inData),
    .io_rightPropDiscard(PEChain_8_io_rightPropDiscard),
    .io_leftOutData(PEChain_8_io_leftOutData),
    .io_rightOutData(PEChain_8_io_rightOutData),
    .io_currDiscard(PEChain_8_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_8_io_toLeftPropDiscard)
  );
  PE_33 PEChain_9 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_9_clock),
    .reset(PEChain_9_reset),
    .io_enableSort(PEChain_9_io_enableSort),
    .io_state(PEChain_9_io_state),
    .io_leftNBR_data(PEChain_9_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_9_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_9_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_9_io_rightNBR_compRes),
    .io_currCell_data(PEChain_9_io_currCell_data),
    .io_currCell_compRes(PEChain_9_io_currCell_compRes),
    .io_lastCell(PEChain_9_io_lastCell),
    .io_active(PEChain_9_io_active),
    .io_discard(PEChain_9_io_discard),
    .io_inData(PEChain_9_io_inData),
    .io_rightPropDiscard(PEChain_9_io_rightPropDiscard),
    .io_leftOutData(PEChain_9_io_leftOutData),
    .io_rightOutData(PEChain_9_io_rightOutData),
    .io_currDiscard(PEChain_9_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_9_io_toLeftPropDiscard)
  );
  PE_34 PEChain_10 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_10_clock),
    .reset(PEChain_10_reset),
    .io_enableSort(PEChain_10_io_enableSort),
    .io_state(PEChain_10_io_state),
    .io_leftNBR_data(PEChain_10_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_10_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_10_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_10_io_rightNBR_compRes),
    .io_currCell_data(PEChain_10_io_currCell_data),
    .io_currCell_compRes(PEChain_10_io_currCell_compRes),
    .io_lastCell(PEChain_10_io_lastCell),
    .io_active(PEChain_10_io_active),
    .io_discard(PEChain_10_io_discard),
    .io_inData(PEChain_10_io_inData),
    .io_rightPropDiscard(PEChain_10_io_rightPropDiscard),
    .io_leftOutData(PEChain_10_io_leftOutData),
    .io_rightOutData(PEChain_10_io_rightOutData),
    .io_currDiscard(PEChain_10_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_10_io_toLeftPropDiscard)
  );
  PE_35 PEChain_11 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_11_clock),
    .reset(PEChain_11_reset),
    .io_enableSort(PEChain_11_io_enableSort),
    .io_state(PEChain_11_io_state),
    .io_leftNBR_data(PEChain_11_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_11_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_11_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_11_io_rightNBR_compRes),
    .io_currCell_data(PEChain_11_io_currCell_data),
    .io_currCell_compRes(PEChain_11_io_currCell_compRes),
    .io_lastCell(PEChain_11_io_lastCell),
    .io_active(PEChain_11_io_active),
    .io_discard(PEChain_11_io_discard),
    .io_inData(PEChain_11_io_inData),
    .io_rightPropDiscard(PEChain_11_io_rightPropDiscard),
    .io_leftOutData(PEChain_11_io_leftOutData),
    .io_rightOutData(PEChain_11_io_rightOutData),
    .io_currDiscard(PEChain_11_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_11_io_toLeftPropDiscard)
  );
  PE_36 PEChain_12 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_12_clock),
    .reset(PEChain_12_reset),
    .io_enableSort(PEChain_12_io_enableSort),
    .io_state(PEChain_12_io_state),
    .io_leftNBR_data(PEChain_12_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_12_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_12_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_12_io_rightNBR_compRes),
    .io_currCell_data(PEChain_12_io_currCell_data),
    .io_currCell_compRes(PEChain_12_io_currCell_compRes),
    .io_lastCell(PEChain_12_io_lastCell),
    .io_active(PEChain_12_io_active),
    .io_discard(PEChain_12_io_discard),
    .io_inData(PEChain_12_io_inData),
    .io_rightPropDiscard(PEChain_12_io_rightPropDiscard),
    .io_leftOutData(PEChain_12_io_leftOutData),
    .io_rightOutData(PEChain_12_io_rightOutData),
    .io_currDiscard(PEChain_12_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_12_io_toLeftPropDiscard)
  );
  PE_37 PEChain_13 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_13_clock),
    .reset(PEChain_13_reset),
    .io_enableSort(PEChain_13_io_enableSort),
    .io_state(PEChain_13_io_state),
    .io_leftNBR_data(PEChain_13_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_13_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_13_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_13_io_rightNBR_compRes),
    .io_currCell_data(PEChain_13_io_currCell_data),
    .io_currCell_compRes(PEChain_13_io_currCell_compRes),
    .io_lastCell(PEChain_13_io_lastCell),
    .io_active(PEChain_13_io_active),
    .io_discard(PEChain_13_io_discard),
    .io_inData(PEChain_13_io_inData),
    .io_rightPropDiscard(PEChain_13_io_rightPropDiscard),
    .io_leftOutData(PEChain_13_io_leftOutData),
    .io_rightOutData(PEChain_13_io_rightOutData),
    .io_currDiscard(PEChain_13_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_13_io_toLeftPropDiscard)
  );
  PE_38 PEChain_14 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_14_clock),
    .reset(PEChain_14_reset),
    .io_enableSort(PEChain_14_io_enableSort),
    .io_state(PEChain_14_io_state),
    .io_leftNBR_data(PEChain_14_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_14_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_14_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_14_io_rightNBR_compRes),
    .io_currCell_data(PEChain_14_io_currCell_data),
    .io_currCell_compRes(PEChain_14_io_currCell_compRes),
    .io_lastCell(PEChain_14_io_lastCell),
    .io_active(PEChain_14_io_active),
    .io_discard(PEChain_14_io_discard),
    .io_inData(PEChain_14_io_inData),
    .io_rightPropDiscard(PEChain_14_io_rightPropDiscard),
    .io_leftOutData(PEChain_14_io_leftOutData),
    .io_rightOutData(PEChain_14_io_rightOutData),
    .io_currDiscard(PEChain_14_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_14_io_toLeftPropDiscard)
  );
  PE_39 PEChain_15 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_15_clock),
    .reset(PEChain_15_reset),
    .io_enableSort(PEChain_15_io_enableSort),
    .io_state(PEChain_15_io_state),
    .io_leftNBR_data(PEChain_15_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_15_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_15_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_15_io_rightNBR_compRes),
    .io_currCell_data(PEChain_15_io_currCell_data),
    .io_currCell_compRes(PEChain_15_io_currCell_compRes),
    .io_lastCell(PEChain_15_io_lastCell),
    .io_active(PEChain_15_io_active),
    .io_discard(PEChain_15_io_discard),
    .io_inData(PEChain_15_io_inData),
    .io_rightPropDiscard(PEChain_15_io_rightPropDiscard),
    .io_leftOutData(PEChain_15_io_leftOutData),
    .io_rightOutData(PEChain_15_io_rightOutData),
    .io_currDiscard(PEChain_15_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_15_io_toLeftPropDiscard)
  );
  PE_40 PEChain_16 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_16_clock),
    .reset(PEChain_16_reset),
    .io_enableSort(PEChain_16_io_enableSort),
    .io_state(PEChain_16_io_state),
    .io_leftNBR_data(PEChain_16_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_16_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_16_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_16_io_rightNBR_compRes),
    .io_currCell_data(PEChain_16_io_currCell_data),
    .io_currCell_compRes(PEChain_16_io_currCell_compRes),
    .io_lastCell(PEChain_16_io_lastCell),
    .io_active(PEChain_16_io_active),
    .io_discard(PEChain_16_io_discard),
    .io_inData(PEChain_16_io_inData),
    .io_rightPropDiscard(PEChain_16_io_rightPropDiscard),
    .io_leftOutData(PEChain_16_io_leftOutData),
    .io_rightOutData(PEChain_16_io_rightOutData),
    .io_currDiscard(PEChain_16_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_16_io_toLeftPropDiscard)
  );
  PE_41 PEChain_17 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_17_clock),
    .reset(PEChain_17_reset),
    .io_enableSort(PEChain_17_io_enableSort),
    .io_state(PEChain_17_io_state),
    .io_leftNBR_data(PEChain_17_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_17_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_17_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_17_io_rightNBR_compRes),
    .io_currCell_data(PEChain_17_io_currCell_data),
    .io_currCell_compRes(PEChain_17_io_currCell_compRes),
    .io_lastCell(PEChain_17_io_lastCell),
    .io_active(PEChain_17_io_active),
    .io_discard(PEChain_17_io_discard),
    .io_inData(PEChain_17_io_inData),
    .io_rightPropDiscard(PEChain_17_io_rightPropDiscard),
    .io_leftOutData(PEChain_17_io_leftOutData),
    .io_rightOutData(PEChain_17_io_rightOutData),
    .io_currDiscard(PEChain_17_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_17_io_toLeftPropDiscard)
  );
  PE_42 PEChain_18 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_18_clock),
    .reset(PEChain_18_reset),
    .io_enableSort(PEChain_18_io_enableSort),
    .io_state(PEChain_18_io_state),
    .io_leftNBR_data(PEChain_18_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_18_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_18_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_18_io_rightNBR_compRes),
    .io_currCell_data(PEChain_18_io_currCell_data),
    .io_currCell_compRes(PEChain_18_io_currCell_compRes),
    .io_lastCell(PEChain_18_io_lastCell),
    .io_active(PEChain_18_io_active),
    .io_discard(PEChain_18_io_discard),
    .io_inData(PEChain_18_io_inData),
    .io_rightPropDiscard(PEChain_18_io_rightPropDiscard),
    .io_leftOutData(PEChain_18_io_leftOutData),
    .io_rightOutData(PEChain_18_io_rightOutData),
    .io_currDiscard(PEChain_18_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_18_io_toLeftPropDiscard)
  );
  PE_43 PEChain_19 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_19_clock),
    .reset(PEChain_19_reset),
    .io_enableSort(PEChain_19_io_enableSort),
    .io_state(PEChain_19_io_state),
    .io_leftNBR_data(PEChain_19_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_19_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_19_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_19_io_rightNBR_compRes),
    .io_currCell_data(PEChain_19_io_currCell_data),
    .io_currCell_compRes(PEChain_19_io_currCell_compRes),
    .io_lastCell(PEChain_19_io_lastCell),
    .io_active(PEChain_19_io_active),
    .io_discard(PEChain_19_io_discard),
    .io_inData(PEChain_19_io_inData),
    .io_rightPropDiscard(PEChain_19_io_rightPropDiscard),
    .io_leftOutData(PEChain_19_io_leftOutData),
    .io_rightOutData(PEChain_19_io_rightOutData),
    .io_currDiscard(PEChain_19_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_19_io_toLeftPropDiscard)
  );
  PE_44 PEChain_20 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_20_clock),
    .reset(PEChain_20_reset),
    .io_enableSort(PEChain_20_io_enableSort),
    .io_state(PEChain_20_io_state),
    .io_leftNBR_data(PEChain_20_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_20_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_20_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_20_io_rightNBR_compRes),
    .io_currCell_data(PEChain_20_io_currCell_data),
    .io_currCell_compRes(PEChain_20_io_currCell_compRes),
    .io_lastCell(PEChain_20_io_lastCell),
    .io_active(PEChain_20_io_active),
    .io_discard(PEChain_20_io_discard),
    .io_inData(PEChain_20_io_inData),
    .io_rightPropDiscard(PEChain_20_io_rightPropDiscard),
    .io_leftOutData(PEChain_20_io_leftOutData),
    .io_rightOutData(PEChain_20_io_rightOutData),
    .io_currDiscard(PEChain_20_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_20_io_toLeftPropDiscard)
  );
  PE_45 PEChain_21 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_21_clock),
    .reset(PEChain_21_reset),
    .io_enableSort(PEChain_21_io_enableSort),
    .io_state(PEChain_21_io_state),
    .io_leftNBR_data(PEChain_21_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_21_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_21_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_21_io_rightNBR_compRes),
    .io_currCell_data(PEChain_21_io_currCell_data),
    .io_currCell_compRes(PEChain_21_io_currCell_compRes),
    .io_lastCell(PEChain_21_io_lastCell),
    .io_active(PEChain_21_io_active),
    .io_discard(PEChain_21_io_discard),
    .io_inData(PEChain_21_io_inData),
    .io_rightPropDiscard(PEChain_21_io_rightPropDiscard),
    .io_leftOutData(PEChain_21_io_leftOutData),
    .io_rightOutData(PEChain_21_io_rightOutData),
    .io_currDiscard(PEChain_21_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_21_io_toLeftPropDiscard)
  );
  PE_46 PEChain_22 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_22_clock),
    .reset(PEChain_22_reset),
    .io_enableSort(PEChain_22_io_enableSort),
    .io_state(PEChain_22_io_state),
    .io_leftNBR_data(PEChain_22_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_22_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_22_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_22_io_rightNBR_compRes),
    .io_currCell_data(PEChain_22_io_currCell_data),
    .io_currCell_compRes(PEChain_22_io_currCell_compRes),
    .io_lastCell(PEChain_22_io_lastCell),
    .io_active(PEChain_22_io_active),
    .io_discard(PEChain_22_io_discard),
    .io_inData(PEChain_22_io_inData),
    .io_rightPropDiscard(PEChain_22_io_rightPropDiscard),
    .io_leftOutData(PEChain_22_io_leftOutData),
    .io_rightOutData(PEChain_22_io_rightOutData),
    .io_currDiscard(PEChain_22_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_22_io_toLeftPropDiscard)
  );
  PE_47 PEChain_23 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_23_clock),
    .reset(PEChain_23_reset),
    .io_enableSort(PEChain_23_io_enableSort),
    .io_state(PEChain_23_io_state),
    .io_leftNBR_data(PEChain_23_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_23_io_leftNBR_compRes),
    .io_currCell_data(PEChain_23_io_currCell_data),
    .io_currCell_compRes(PEChain_23_io_currCell_compRes),
    .io_lastCell(PEChain_23_io_lastCell),
    .io_active(PEChain_23_io_active),
    .io_discard(PEChain_23_io_discard),
    .io_inData(PEChain_23_io_inData),
    .io_leftOutData(PEChain_23_io_leftOutData),
    .io_currDiscard(PEChain_23_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_23_io_toLeftPropDiscard)
  );
  assign _T_1 = lisSizeReg - 6'h1; // @[LinearSorter.scala 86:43]
  assign _T_96 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_98 = cntInData + 5'h1; // @[LinearSorter.scala 92:28]
  assign _T_99 = state == 2'h0; // @[LinearSorter.scala 94:20]
  assign _GEN_111 = {{1'd0}, cntInData}; // @[LinearSorter.scala 98:19]
  assign _T_102 = _GEN_111 == _T_1; // @[LinearSorter.scala 98:19]
  assign _T_104 = _T_102 & _T_96; // @[LinearSorter.scala 98:42]
  assign _T_113 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_7 = _T_96 ? 2'h1 : state; // @[LinearSorter.scala 117:27]
  assign _T_115 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign fireLastIn = io_lastIn & _T_96; // @[LinearSorter.scala 111:30]
  assign _GEN_8 = fireLastIn ? 2'h2 : state; // @[LinearSorter.scala 120:62]
  assign _T_117 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_112 = {{1'd0}, cntOutData}; // @[LinearSorter.scala 125:28]
  assign _T_120 = _GEN_112 == _T_1; // @[LinearSorter.scala 125:28]
  assign _GEN_9 = _T_120 ? 2'h0 : state; // @[LinearSorter.scala 125:50]
  assign _GEN_10 = _T_117 ? _GEN_9 : state; // @[Conditional.scala 39:67]
  assign _GEN_11 = _T_115 ? _GEN_8 : _GEN_10; // @[Conditional.scala 39:67]
  assign state_next = _T_113 ? _GEN_7 : _GEN_11; // @[Conditional.scala 40:58]
  assign _T_105 = state_next == 2'h0; // @[LinearSorter.scala 101:25]
  assign _GEN_2 = _T_105 ? 1'h0 : initialInDone; // @[LinearSorter.scala 101:36]
  assign _GEN_3 = _T_104 | _GEN_2; // @[LinearSorter.scala 98:59]
  assign _T_106 = io_out_valid & io_out_ready; // @[LinearSorter.scala 106:29]
  assign _T_107 = state == 2'h2; // @[LinearSorter.scala 106:54]
  assign enable = _T_106 & _T_107; // @[LinearSorter.scala 106:45]
  assign _T_109 = cntOutData == 5'h17; // @[LISutil.scala 13:24]
  assign _T_111 = cntOutData + 5'h1; // @[LISutil.scala 14:22]
  assign _T_121 = state_next != 2'h2; // @[LinearSorter.scala 137:33]
  assign outputData_0 = PEChain_0_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign outputData_1 = PEChain_1_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_16 = 5'h1 == _T_1[4:0] ? $signed(outputData_1) : $signed(outputData_0); // @[LinearSorter.scala 137:21]
  assign outputData_2 = PEChain_2_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_17 = 5'h2 == _T_1[4:0] ? $signed(outputData_2) : $signed(_GEN_16); // @[LinearSorter.scala 137:21]
  assign outputData_3 = PEChain_3_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_18 = 5'h3 == _T_1[4:0] ? $signed(outputData_3) : $signed(_GEN_17); // @[LinearSorter.scala 137:21]
  assign outputData_4 = PEChain_4_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_19 = 5'h4 == _T_1[4:0] ? $signed(outputData_4) : $signed(_GEN_18); // @[LinearSorter.scala 137:21]
  assign outputData_5 = PEChain_5_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_20 = 5'h5 == _T_1[4:0] ? $signed(outputData_5) : $signed(_GEN_19); // @[LinearSorter.scala 137:21]
  assign outputData_6 = PEChain_6_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_21 = 5'h6 == _T_1[4:0] ? $signed(outputData_6) : $signed(_GEN_20); // @[LinearSorter.scala 137:21]
  assign outputData_7 = PEChain_7_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_22 = 5'h7 == _T_1[4:0] ? $signed(outputData_7) : $signed(_GEN_21); // @[LinearSorter.scala 137:21]
  assign outputData_8 = PEChain_8_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_23 = 5'h8 == _T_1[4:0] ? $signed(outputData_8) : $signed(_GEN_22); // @[LinearSorter.scala 137:21]
  assign outputData_9 = PEChain_9_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_24 = 5'h9 == _T_1[4:0] ? $signed(outputData_9) : $signed(_GEN_23); // @[LinearSorter.scala 137:21]
  assign outputData_10 = PEChain_10_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_25 = 5'ha == _T_1[4:0] ? $signed(outputData_10) : $signed(_GEN_24); // @[LinearSorter.scala 137:21]
  assign outputData_11 = PEChain_11_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_26 = 5'hb == _T_1[4:0] ? $signed(outputData_11) : $signed(_GEN_25); // @[LinearSorter.scala 137:21]
  assign outputData_12 = PEChain_12_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_27 = 5'hc == _T_1[4:0] ? $signed(outputData_12) : $signed(_GEN_26); // @[LinearSorter.scala 137:21]
  assign outputData_13 = PEChain_13_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_28 = 5'hd == _T_1[4:0] ? $signed(outputData_13) : $signed(_GEN_27); // @[LinearSorter.scala 137:21]
  assign outputData_14 = PEChain_14_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_29 = 5'he == _T_1[4:0] ? $signed(outputData_14) : $signed(_GEN_28); // @[LinearSorter.scala 137:21]
  assign outputData_15 = PEChain_15_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_30 = 5'hf == _T_1[4:0] ? $signed(outputData_15) : $signed(_GEN_29); // @[LinearSorter.scala 137:21]
  assign outputData_16 = PEChain_16_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_31 = 5'h10 == _T_1[4:0] ? $signed(outputData_16) : $signed(_GEN_30); // @[LinearSorter.scala 137:21]
  assign outputData_17 = PEChain_17_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_32 = 5'h11 == _T_1[4:0] ? $signed(outputData_17) : $signed(_GEN_31); // @[LinearSorter.scala 137:21]
  assign outputData_18 = PEChain_18_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_33 = 5'h12 == _T_1[4:0] ? $signed(outputData_18) : $signed(_GEN_32); // @[LinearSorter.scala 137:21]
  assign outputData_19 = PEChain_19_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_34 = 5'h13 == _T_1[4:0] ? $signed(outputData_19) : $signed(_GEN_33); // @[LinearSorter.scala 137:21]
  assign outputData_20 = PEChain_20_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_35 = 5'h14 == _T_1[4:0] ? $signed(outputData_20) : $signed(_GEN_34); // @[LinearSorter.scala 137:21]
  assign outputData_21 = PEChain_21_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_36 = 5'h15 == _T_1[4:0] ? $signed(outputData_21) : $signed(_GEN_35); // @[LinearSorter.scala 137:21]
  assign outputData_22 = PEChain_22_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_37 = 5'h16 == _T_1[4:0] ? $signed(outputData_22) : $signed(_GEN_36); // @[LinearSorter.scala 137:21]
  assign outputData_23 = PEChain_23_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_38 = 5'h17 == _T_1[4:0] ? $signed(outputData_23) : $signed(_GEN_37); // @[LinearSorter.scala 137:21]
  assign _T_132 = 5'h0 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_39 = _T_132 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_136 = _T_107 & io_out_ready; // @[LinearSorter.scala 168:63]
  assign _T_142 = 5'h1 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_41 = _T_142 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_152 = 5'h2 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_43 = _T_152 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_162 = 5'h3 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_45 = _T_162 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_172 = 5'h4 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_47 = _T_172 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_182 = 5'h5 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_49 = _T_182 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_192 = 5'h6 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_51 = _T_192 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_202 = 5'h7 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_53 = _T_202 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_212 = 5'h8 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_55 = _T_212 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_222 = 5'h9 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_57 = _T_222 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_232 = 5'ha == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_59 = _T_232 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_242 = 5'hb == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_61 = _T_242 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_252 = 5'hc == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_63 = _T_252 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_262 = 5'hd == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_65 = _T_262 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_272 = 5'he == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_67 = _T_272 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_282 = 5'hf == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_69 = _T_282 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_292 = 5'h10 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_71 = _T_292 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_302 = 5'h11 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_73 = _T_302 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_312 = 5'h12 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_75 = _T_312 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_322 = 5'h13 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_77 = _T_322 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_332 = 5'h14 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_79 = _T_332 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_342 = 5'h15 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_81 = _T_342 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_352 = 5'h16 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_83 = _T_352 & initialInDone; // @[LinearSorter.scala 160:80]
  assign _T_362 = 5'h17 == io_discardPos; // @[LinearSorter.scala 160:26]
  assign _GEN_85 = _T_362 & initialInDone; // @[LinearSorter.scala 160:80]
  assign discardSignals_2 = PEChain_2_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_1 = PEChain_1_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_0 = PEChain_0_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_5 = PEChain_5_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_4 = PEChain_4_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_3 = PEChain_3_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_372 = {discardSignals_5,discardSignals_4,discardSignals_3,discardSignals_2,discardSignals_1,discardSignals_0}; // @[LinearSorter.scala 177:50]
  assign discardSignals_8 = PEChain_8_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_7 = PEChain_7_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_6 = PEChain_6_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_11 = PEChain_11_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_10 = PEChain_10_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_9 = PEChain_9_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_378 = {discardSignals_11,discardSignals_10,discardSignals_9,discardSignals_8,discardSignals_7,discardSignals_6,_T_372}; // @[LinearSorter.scala 177:50]
  assign discardSignals_14 = PEChain_14_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_13 = PEChain_13_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_12 = PEChain_12_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_17 = PEChain_17_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_16 = PEChain_16_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_15 = PEChain_15_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_383 = {discardSignals_17,discardSignals_16,discardSignals_15,discardSignals_14,discardSignals_13,discardSignals_12}; // @[LinearSorter.scala 177:50]
  assign discardSignals_20 = PEChain_20_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_19 = PEChain_19_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_18 = PEChain_18_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_23 = PEChain_23_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_22 = PEChain_22_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_21 = PEChain_21_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_390 = {discardSignals_23,discardSignals_22,discardSignals_21,discardSignals_20,discardSignals_19,discardSignals_18,_T_383,_T_378}; // @[LinearSorter.scala 177:50]
  assign _T_415 = _T_390[22] ? 5'h16 : 5'h17; // @[Mux.scala 47:69]
  assign _T_416 = _T_390[21] ? 5'h15 : _T_415; // @[Mux.scala 47:69]
  assign _T_417 = _T_390[20] ? 5'h14 : _T_416; // @[Mux.scala 47:69]
  assign _T_418 = _T_390[19] ? 5'h13 : _T_417; // @[Mux.scala 47:69]
  assign _T_419 = _T_390[18] ? 5'h12 : _T_418; // @[Mux.scala 47:69]
  assign _T_420 = _T_390[17] ? 5'h11 : _T_419; // @[Mux.scala 47:69]
  assign _T_421 = _T_390[16] ? 5'h10 : _T_420; // @[Mux.scala 47:69]
  assign _T_422 = _T_390[15] ? 5'hf : _T_421; // @[Mux.scala 47:69]
  assign _T_423 = _T_390[14] ? 5'he : _T_422; // @[Mux.scala 47:69]
  assign _T_424 = _T_390[13] ? 5'hd : _T_423; // @[Mux.scala 47:69]
  assign _T_425 = _T_390[12] ? 5'hc : _T_424; // @[Mux.scala 47:69]
  assign _T_426 = _T_390[11] ? 5'hb : _T_425; // @[Mux.scala 47:69]
  assign _T_427 = _T_390[10] ? 5'ha : _T_426; // @[Mux.scala 47:69]
  assign _T_428 = _T_390[9] ? 5'h9 : _T_427; // @[Mux.scala 47:69]
  assign _T_429 = _T_390[8] ? 5'h8 : _T_428; // @[Mux.scala 47:69]
  assign _T_430 = _T_390[7] ? 5'h7 : _T_429; // @[Mux.scala 47:69]
  assign _T_431 = _T_390[6] ? 5'h6 : _T_430; // @[Mux.scala 47:69]
  assign _T_432 = _T_390[5] ? 5'h5 : _T_431; // @[Mux.scala 47:69]
  assign _T_433 = _T_390[4] ? 5'h4 : _T_432; // @[Mux.scala 47:69]
  assign _T_434 = _T_390[3] ? 5'h3 : _T_433; // @[Mux.scala 47:69]
  assign _T_435 = _T_390[2] ? 5'h2 : _T_434; // @[Mux.scala 47:69]
  assign _T_436 = _T_390[1] ? 5'h1 : _T_435; // @[Mux.scala 47:69]
  assign getDiscarded = _T_390[0] ? 5'h0 : _T_436; // @[Mux.scala 47:69]
  assign _T_438 = state != 2'h2; // @[LinearSorter.scala 199:49]
  assign _GEN_88 = 5'h1 == getDiscarded ? $signed(outputData_1) : $signed(outputData_0); // @[LinearSorter.scala 206:15]
  assign _GEN_89 = 5'h2 == getDiscarded ? $signed(outputData_2) : $signed(_GEN_88); // @[LinearSorter.scala 206:15]
  assign _GEN_90 = 5'h3 == getDiscarded ? $signed(outputData_3) : $signed(_GEN_89); // @[LinearSorter.scala 206:15]
  assign _GEN_91 = 5'h4 == getDiscarded ? $signed(outputData_4) : $signed(_GEN_90); // @[LinearSorter.scala 206:15]
  assign _GEN_92 = 5'h5 == getDiscarded ? $signed(outputData_5) : $signed(_GEN_91); // @[LinearSorter.scala 206:15]
  assign _GEN_93 = 5'h6 == getDiscarded ? $signed(outputData_6) : $signed(_GEN_92); // @[LinearSorter.scala 206:15]
  assign _GEN_94 = 5'h7 == getDiscarded ? $signed(outputData_7) : $signed(_GEN_93); // @[LinearSorter.scala 206:15]
  assign _GEN_95 = 5'h8 == getDiscarded ? $signed(outputData_8) : $signed(_GEN_94); // @[LinearSorter.scala 206:15]
  assign _GEN_96 = 5'h9 == getDiscarded ? $signed(outputData_9) : $signed(_GEN_95); // @[LinearSorter.scala 206:15]
  assign _GEN_97 = 5'ha == getDiscarded ? $signed(outputData_10) : $signed(_GEN_96); // @[LinearSorter.scala 206:15]
  assign _GEN_98 = 5'hb == getDiscarded ? $signed(outputData_11) : $signed(_GEN_97); // @[LinearSorter.scala 206:15]
  assign _GEN_99 = 5'hc == getDiscarded ? $signed(outputData_12) : $signed(_GEN_98); // @[LinearSorter.scala 206:15]
  assign _GEN_100 = 5'hd == getDiscarded ? $signed(outputData_13) : $signed(_GEN_99); // @[LinearSorter.scala 206:15]
  assign _GEN_101 = 5'he == getDiscarded ? $signed(outputData_14) : $signed(_GEN_100); // @[LinearSorter.scala 206:15]
  assign _GEN_102 = 5'hf == getDiscarded ? $signed(outputData_15) : $signed(_GEN_101); // @[LinearSorter.scala 206:15]
  assign _GEN_103 = 5'h10 == getDiscarded ? $signed(outputData_16) : $signed(_GEN_102); // @[LinearSorter.scala 206:15]
  assign _GEN_104 = 5'h11 == getDiscarded ? $signed(outputData_17) : $signed(_GEN_103); // @[LinearSorter.scala 206:15]
  assign _GEN_105 = 5'h12 == getDiscarded ? $signed(outputData_18) : $signed(_GEN_104); // @[LinearSorter.scala 206:15]
  assign _GEN_106 = 5'h13 == getDiscarded ? $signed(outputData_19) : $signed(_GEN_105); // @[LinearSorter.scala 206:15]
  assign _GEN_107 = 5'h14 == getDiscarded ? $signed(outputData_20) : $signed(_GEN_106); // @[LinearSorter.scala 206:15]
  assign _GEN_108 = 5'h15 == getDiscarded ? $signed(outputData_21) : $signed(_GEN_107); // @[LinearSorter.scala 206:15]
  assign _GEN_109 = 5'h16 == getDiscarded ? $signed(outputData_22) : $signed(_GEN_108); // @[LinearSorter.scala 206:15]
  assign _T_444 = ~initialInDone; // @[LinearSorter.scala 208:18]
  assign _T_446 = io_out_ready & _T_438; // @[LinearSorter.scala 208:49]
  assign _T_448 = initialInDone & io_in_valid; // @[LinearSorter.scala 209:33]
  assign io_in_ready = _T_444 | _T_446; // @[LinearSorter.scala 208:15]
  assign io_out_valid = _T_448 | _T_107; // @[LinearSorter.scala 209:16]
  assign io_out_bits = 5'h17 == getDiscarded ? $signed(outputData_23) : $signed(_GEN_109); // @[LinearSorter.scala 206:15]
  assign io_lastOut = _GEN_112 == _T_1; // @[LinearSorter.scala 207:15]
  assign io_sortedData_0 = PEChain_0_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_1 = PEChain_1_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_2 = PEChain_2_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_3 = PEChain_3_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_4 = PEChain_4_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_5 = PEChain_5_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_6 = PEChain_6_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_7 = PEChain_7_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_8 = PEChain_8_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_9 = PEChain_9_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_10 = PEChain_10_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_11 = PEChain_11_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_12 = PEChain_12_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_13 = PEChain_13_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_14 = PEChain_14_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_15 = PEChain_15_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_16 = PEChain_16_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_17 = PEChain_17_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_18 = PEChain_18_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_19 = PEChain_19_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_20 = PEChain_20_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_21 = PEChain_21_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_22 = PEChain_22_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_23 = PEChain_23_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sorterFull = initialInDone & _T_438; // @[LinearSorter.scala 199:23]
  assign io_sorterEmpty = state == 2'h0; // @[LinearSorter.scala 202:24]
  assign PEChain_0_clock = clock;
  assign PEChain_0_reset = reset;
  assign PEChain_0_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_0_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_0_io_rightNBR_data = PEChain_1_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_0_io_rightNBR_compRes = PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_0_io_lastCell = 6'h0 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_0_io_discard = _T_107 ? initialInDone : _GEN_39; // @[LinearSorter.scala 156:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_0_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_0_io_rightPropDiscard = PEChain_1_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_1_clock = clock;
  assign PEChain_1_reset = reset;
  assign PEChain_1_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_1_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_1_io_leftNBR_data = PEChain_0_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_1_io_leftNBR_compRes = PEChain_0_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_1_io_rightNBR_data = PEChain_2_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_1_io_rightNBR_compRes = PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_1_io_lastCell = 6'h1 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_1_io_active = 6'h1 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_1_io_discard = _T_107 ? 1'h0 : _GEN_41; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_1_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_1_io_rightPropDiscard = PEChain_2_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_2_clock = clock;
  assign PEChain_2_reset = reset;
  assign PEChain_2_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_2_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_2_io_leftNBR_data = PEChain_1_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_2_io_leftNBR_compRes = PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_2_io_rightNBR_data = PEChain_3_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_2_io_rightNBR_compRes = PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_2_io_lastCell = 6'h2 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_2_io_active = 6'h2 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_2_io_discard = _T_107 ? 1'h0 : _GEN_43; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_2_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_2_io_rightPropDiscard = PEChain_3_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_3_clock = clock;
  assign PEChain_3_reset = reset;
  assign PEChain_3_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_3_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_3_io_leftNBR_data = PEChain_2_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_3_io_leftNBR_compRes = PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_3_io_rightNBR_data = PEChain_4_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_3_io_rightNBR_compRes = PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_3_io_lastCell = 6'h3 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_3_io_active = 6'h3 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_3_io_discard = _T_107 ? 1'h0 : _GEN_45; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_3_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_3_io_rightPropDiscard = PEChain_4_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_4_clock = clock;
  assign PEChain_4_reset = reset;
  assign PEChain_4_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_4_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_4_io_leftNBR_data = PEChain_3_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_4_io_leftNBR_compRes = PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_4_io_rightNBR_data = PEChain_5_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_4_io_rightNBR_compRes = PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_4_io_lastCell = 6'h4 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_4_io_active = 6'h4 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_4_io_discard = _T_107 ? 1'h0 : _GEN_47; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_4_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_4_io_rightPropDiscard = PEChain_5_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_5_clock = clock;
  assign PEChain_5_reset = reset;
  assign PEChain_5_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_5_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_5_io_leftNBR_data = PEChain_4_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_5_io_leftNBR_compRes = PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_5_io_rightNBR_data = PEChain_6_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_5_io_rightNBR_compRes = PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_5_io_lastCell = 6'h5 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_5_io_active = 6'h5 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_5_io_discard = _T_107 ? 1'h0 : _GEN_49; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_5_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_5_io_rightPropDiscard = PEChain_6_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_6_clock = clock;
  assign PEChain_6_reset = reset;
  assign PEChain_6_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_6_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_6_io_leftNBR_data = PEChain_5_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_6_io_leftNBR_compRes = PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_6_io_rightNBR_data = PEChain_7_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_6_io_rightNBR_compRes = PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_6_io_lastCell = 6'h6 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_6_io_active = 6'h6 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_6_io_discard = _T_107 ? 1'h0 : _GEN_51; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_6_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_6_io_rightPropDiscard = PEChain_7_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_7_clock = clock;
  assign PEChain_7_reset = reset;
  assign PEChain_7_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_7_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_7_io_leftNBR_data = PEChain_6_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_7_io_leftNBR_compRes = PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_7_io_rightNBR_data = PEChain_8_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_7_io_rightNBR_compRes = PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_7_io_lastCell = 6'h7 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_7_io_active = 6'h7 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_7_io_discard = _T_107 ? 1'h0 : _GEN_53; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_7_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_7_io_rightPropDiscard = PEChain_8_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_8_clock = clock;
  assign PEChain_8_reset = reset;
  assign PEChain_8_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_8_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_8_io_leftNBR_data = PEChain_7_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_8_io_leftNBR_compRes = PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_8_io_rightNBR_data = PEChain_9_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_8_io_rightNBR_compRes = PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_8_io_lastCell = 6'h8 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_8_io_active = 6'h8 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_8_io_discard = _T_107 ? 1'h0 : _GEN_55; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_8_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_8_io_rightPropDiscard = PEChain_9_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_9_clock = clock;
  assign PEChain_9_reset = reset;
  assign PEChain_9_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_9_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_9_io_leftNBR_data = PEChain_8_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_9_io_leftNBR_compRes = PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_9_io_rightNBR_data = PEChain_10_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_9_io_rightNBR_compRes = PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_9_io_lastCell = 6'h9 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_9_io_active = 6'h9 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_9_io_discard = _T_107 ? 1'h0 : _GEN_57; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_9_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_9_io_rightPropDiscard = PEChain_10_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_10_clock = clock;
  assign PEChain_10_reset = reset;
  assign PEChain_10_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_10_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_10_io_leftNBR_data = PEChain_9_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_10_io_leftNBR_compRes = PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_10_io_rightNBR_data = PEChain_11_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_10_io_rightNBR_compRes = PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_10_io_lastCell = 6'ha == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_10_io_active = 6'ha <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_10_io_discard = _T_107 ? 1'h0 : _GEN_59; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_10_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_10_io_rightPropDiscard = PEChain_11_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_11_clock = clock;
  assign PEChain_11_reset = reset;
  assign PEChain_11_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_11_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_11_io_leftNBR_data = PEChain_10_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_11_io_leftNBR_compRes = PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_11_io_rightNBR_data = PEChain_12_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_11_io_rightNBR_compRes = PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_11_io_lastCell = 6'hb == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_11_io_active = 6'hb <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_11_io_discard = _T_107 ? 1'h0 : _GEN_61; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_11_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_11_io_rightPropDiscard = PEChain_12_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_12_clock = clock;
  assign PEChain_12_reset = reset;
  assign PEChain_12_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_12_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_12_io_leftNBR_data = PEChain_11_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_12_io_leftNBR_compRes = PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_12_io_rightNBR_data = PEChain_13_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_12_io_rightNBR_compRes = PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_12_io_lastCell = 6'hc == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_12_io_active = 6'hc <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_12_io_discard = _T_107 ? 1'h0 : _GEN_63; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_12_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_12_io_rightPropDiscard = PEChain_13_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_13_clock = clock;
  assign PEChain_13_reset = reset;
  assign PEChain_13_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_13_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_13_io_leftNBR_data = PEChain_12_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_13_io_leftNBR_compRes = PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_13_io_rightNBR_data = PEChain_14_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_13_io_rightNBR_compRes = PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_13_io_lastCell = 6'hd == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_13_io_active = 6'hd <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_13_io_discard = _T_107 ? 1'h0 : _GEN_65; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_13_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_13_io_rightPropDiscard = PEChain_14_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_14_clock = clock;
  assign PEChain_14_reset = reset;
  assign PEChain_14_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_14_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_14_io_leftNBR_data = PEChain_13_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_14_io_leftNBR_compRes = PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_14_io_rightNBR_data = PEChain_15_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_14_io_rightNBR_compRes = PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_14_io_lastCell = 6'he == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_14_io_active = 6'he <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_14_io_discard = _T_107 ? 1'h0 : _GEN_67; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_14_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_14_io_rightPropDiscard = PEChain_15_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_15_clock = clock;
  assign PEChain_15_reset = reset;
  assign PEChain_15_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_15_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_15_io_leftNBR_data = PEChain_14_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_15_io_leftNBR_compRes = PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_15_io_rightNBR_data = PEChain_16_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_15_io_rightNBR_compRes = PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_15_io_lastCell = 6'hf == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_15_io_active = 6'hf <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_15_io_discard = _T_107 ? 1'h0 : _GEN_69; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_15_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_15_io_rightPropDiscard = PEChain_16_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_16_clock = clock;
  assign PEChain_16_reset = reset;
  assign PEChain_16_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_16_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_16_io_leftNBR_data = PEChain_15_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_16_io_leftNBR_compRes = PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_16_io_rightNBR_data = PEChain_17_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_16_io_rightNBR_compRes = PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_16_io_lastCell = 6'h10 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_16_io_active = 6'h10 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_16_io_discard = _T_107 ? 1'h0 : _GEN_71; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_16_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_16_io_rightPropDiscard = PEChain_17_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_17_clock = clock;
  assign PEChain_17_reset = reset;
  assign PEChain_17_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_17_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_17_io_leftNBR_data = PEChain_16_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_17_io_leftNBR_compRes = PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_17_io_rightNBR_data = PEChain_18_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_17_io_rightNBR_compRes = PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_17_io_lastCell = 6'h11 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_17_io_active = 6'h11 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_17_io_discard = _T_107 ? 1'h0 : _GEN_73; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_17_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_17_io_rightPropDiscard = PEChain_18_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_18_clock = clock;
  assign PEChain_18_reset = reset;
  assign PEChain_18_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_18_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_18_io_leftNBR_data = PEChain_17_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_18_io_leftNBR_compRes = PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_18_io_rightNBR_data = PEChain_19_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_18_io_rightNBR_compRes = PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_18_io_lastCell = 6'h12 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_18_io_active = 6'h12 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_18_io_discard = _T_107 ? 1'h0 : _GEN_75; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_18_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_18_io_rightPropDiscard = PEChain_19_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_19_clock = clock;
  assign PEChain_19_reset = reset;
  assign PEChain_19_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_19_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_19_io_leftNBR_data = PEChain_18_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_19_io_leftNBR_compRes = PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_19_io_rightNBR_data = PEChain_20_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_19_io_rightNBR_compRes = PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_19_io_lastCell = 6'h13 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_19_io_active = 6'h13 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_19_io_discard = _T_107 ? 1'h0 : _GEN_77; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_19_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_19_io_rightPropDiscard = PEChain_20_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_20_clock = clock;
  assign PEChain_20_reset = reset;
  assign PEChain_20_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_20_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_20_io_leftNBR_data = PEChain_19_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_20_io_leftNBR_compRes = PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_20_io_rightNBR_data = PEChain_21_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_20_io_rightNBR_compRes = PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_20_io_lastCell = 6'h14 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_20_io_active = 6'h14 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_20_io_discard = _T_107 ? 1'h0 : _GEN_79; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_20_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_20_io_rightPropDiscard = PEChain_21_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_21_clock = clock;
  assign PEChain_21_reset = reset;
  assign PEChain_21_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_21_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_21_io_leftNBR_data = PEChain_20_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_21_io_leftNBR_compRes = PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_21_io_rightNBR_data = PEChain_22_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_21_io_rightNBR_compRes = PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_21_io_lastCell = 6'h15 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_21_io_active = 6'h15 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_21_io_discard = _T_107 ? 1'h0 : _GEN_81; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_21_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_21_io_rightPropDiscard = PEChain_22_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_22_clock = clock;
  assign PEChain_22_reset = reset;
  assign PEChain_22_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_22_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_22_io_leftNBR_data = PEChain_21_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_22_io_leftNBR_compRes = PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_22_io_rightNBR_data = PEChain_23_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_22_io_rightNBR_compRes = PEChain_23_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_22_io_lastCell = 6'h16 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_22_io_active = 6'h16 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_22_io_discard = _T_107 ? 1'h0 : _GEN_83; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_22_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_22_io_rightPropDiscard = PEChain_23_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_23_clock = clock;
  assign PEChain_23_reset = reset;
  assign PEChain_23_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_23_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_23_io_leftNBR_data = PEChain_22_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_23_io_leftNBR_compRes = PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_23_io_lastCell = 6'h17 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_23_io_active = 6'h17 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_23_io_discard = _T_107 ? 1'h0 : _GEN_85; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_23_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntInData = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  lisSizeReg = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cntOutData = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_3;
    end
    if (reset) begin
      cntInData <= 5'h0;
    end else if (_T_96) begin
      cntInData <= _T_98;
    end else if (_T_99) begin
      cntInData <= 5'h0;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_113) begin
      if (_T_96) begin
        state <= 2'h1;
      end
    end else if (_T_115) begin
      if (fireLastIn) begin
        state <= 2'h2;
      end
    end else if (_T_117) begin
      if (_T_120) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      lisSizeReg <= 6'h18;
    end else if (_T_113) begin
      lisSizeReg <= io_lisSize;
    end
    if (reset) begin
      cntOutData <= 5'h0;
    end else if (_T_99) begin
      cntOutData <= 5'h0;
    end else if (enable) begin
      if (_T_109) begin
        cntOutData <= 5'h0;
      end else begin
        cntOutData <= _T_111;
      end
    end
  end
endmodule
module AXI4LISBlock_1(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  lis_clock; // @[LISDspBlock.scala 55:21]
  wire  lis_reset; // @[LISDspBlock.scala 55:21]
  wire  lis_io_in_ready; // @[LISDspBlock.scala 55:21]
  wire  lis_io_in_valid; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_in_bits; // @[LISDspBlock.scala 55:21]
  wire  lis_io_lastIn; // @[LISDspBlock.scala 55:21]
  wire  lis_io_out_ready; // @[LISDspBlock.scala 55:21]
  wire  lis_io_out_valid; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_out_bits; // @[LISDspBlock.scala 55:21]
  wire  lis_io_lastOut; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_0; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_1; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_2; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_3; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_4; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_5; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_6; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_7; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_8; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_9; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_10; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_11; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_12; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_13; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_14; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_15; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_16; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_17; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_18; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_19; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_20; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_21; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_22; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_23; // @[LISDspBlock.scala 55:21]
  wire  lis_io_sorterFull; // @[LISDspBlock.scala 55:21]
  wire  lis_io_sorterEmpty; // @[LISDspBlock.scala 55:21]
  wire [5:0] lis_io_lisSize; // @[LISDspBlock.scala 55:21]
  wire [4:0] lis_io_discardPos; // @[LISDspBlock.scala 55:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  sortDir; // @[LISDspBlock.scala 58:26]
  reg [31:0] _RAND_0;
  reg  flushData; // @[LISDspBlock.scala 59:28]
  reg [31:0] _RAND_1;
  reg [4:0] discardPos; // @[LISDspBlock.scala 60:29]
  reg [31:0] _RAND_2;
  reg [4:0] sendOnOutput; // @[LISDspBlock.scala 61:31]
  reg [31:0] _RAND_3;
  reg [4:0] lisSize; // @[LISDspBlock.scala 62:26]
  reg [31:0] _RAND_4;
  reg  sorterFull; // @[LISDspBlock.scala 65:29]
  reg [31:0] _RAND_5;
  reg  sorterEmpty; // @[LISDspBlock.scala 66:30]
  reg [31:0] _RAND_6;
  wire [31:0] _T_2; // @[LISDspBlock.scala 71:44]
  wire [15:0] _GEN_0; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_1; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_2; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_3; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_4; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_5; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_6; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_7; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_8; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_9; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_10; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_11; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_12; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_13; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_14; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_15; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_16; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_17; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_18; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_19; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_20; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_21; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_22; // @[LISDspBlock.scala 92:82]
  wire [15:0] _T_4; // @[LISDspBlock.scala 92:82]
  wire  _T_7; // @[RegisterRouter.scala 40:39]
  wire  _T_8; // @[RegisterRouter.scala 40:26]
  wire  _T_9; // @[RegisterRouter.scala 42:29]
  wire  _T_52_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_16; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_281; // @[Cat.scala 29:58]
  wire [5:0] _T_56; // @[RegisterRouter.scala 59:16]
  wire  _T_64; // @[RegisterRouter.scala 59:16]
  wire  _T_10; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_19; // @[OneHot.scala 65:12]
  wire [1:0] _T_21; // @[Misc.scala 200:81]
  wire  _T_22; // @[Misc.scala 204:21]
  wire  _T_25; // @[Misc.scala 209:20]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_30; // @[Misc.scala 213:38]
  wire  _T_31; // @[Misc.scala 213:29]
  wire  _T_34; // @[Misc.scala 209:20]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 212:27]
  wire  _T_45; // @[Misc.scala 213:38]
  wire  _T_46; // @[Misc.scala 213:29]
  wire [3:0] _T_49; // @[Cat.scala 29:58]
  wire [3:0] _T_51; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_300; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_282; // @[OneHot.scala 58:35]
  wire  _T_347; // @[RegisterRouter.scala 59:16]
  wire  _T_349; // @[RegisterRouter.scala 59:16]
  wire  _T_350; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _GEN_24; // @[RegField.scala 134:88]
  wire  _T_154; // @[RegisterRouter.scala 59:16]
  wire  _T_354; // @[RegisterRouter.scala 59:16]
  wire  _T_355; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire  _T_359; // @[RegisterRouter.scala 59:16]
  wire  _T_360; // @[RegisterRouter.scala 59:16]
  wire  _T_207; // @[RegisterRouter.scala 59:16]
  wire  _T_364; // @[RegisterRouter.scala 59:16]
  wire  _T_365; // @[RegisterRouter.scala 59:16]
  wire  _T_230; // @[RegisterRouter.scala 59:16]
  wire  _T_369; // @[RegisterRouter.scala 59:16]
  wire  _T_370; // @[RegisterRouter.scala 59:16]
  wire  _T_253; // @[RegisterRouter.scala 59:16]
  wire  _GEN_62; // @[MuxLiteral.scala 48:10]
  wire  _GEN_63; // @[MuxLiteral.scala 48:10]
  wire  _GEN_64; // @[MuxLiteral.scala 48:10]
  wire  _GEN_65; // @[MuxLiteral.scala 48:10]
  wire  _GEN_66; // @[MuxLiteral.scala 48:10]
  wire  _GEN_67; // @[MuxLiteral.scala 48:10]
  wire  _GEN_77; // @[MuxLiteral.scala 48:10]
  wire  _GEN_68; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_70; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_71; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_72; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_73; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_74; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_75; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_76; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_494; // @[RegisterRouter.scala 59:16]
  wire  _T_495_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_495_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_498; // @[RegisterRouter.scala 65:29]
  LinearSorter_1 lis ( // @[LISDspBlock.scala 55:21]
    .clock(lis_clock),
    .reset(lis_reset),
    .io_in_ready(lis_io_in_ready),
    .io_in_valid(lis_io_in_valid),
    .io_in_bits(lis_io_in_bits),
    .io_lastIn(lis_io_lastIn),
    .io_out_ready(lis_io_out_ready),
    .io_out_valid(lis_io_out_valid),
    .io_out_bits(lis_io_out_bits),
    .io_lastOut(lis_io_lastOut),
    .io_sortedData_0(lis_io_sortedData_0),
    .io_sortedData_1(lis_io_sortedData_1),
    .io_sortedData_2(lis_io_sortedData_2),
    .io_sortedData_3(lis_io_sortedData_3),
    .io_sortedData_4(lis_io_sortedData_4),
    .io_sortedData_5(lis_io_sortedData_5),
    .io_sortedData_6(lis_io_sortedData_6),
    .io_sortedData_7(lis_io_sortedData_7),
    .io_sortedData_8(lis_io_sortedData_8),
    .io_sortedData_9(lis_io_sortedData_9),
    .io_sortedData_10(lis_io_sortedData_10),
    .io_sortedData_11(lis_io_sortedData_11),
    .io_sortedData_12(lis_io_sortedData_12),
    .io_sortedData_13(lis_io_sortedData_13),
    .io_sortedData_14(lis_io_sortedData_14),
    .io_sortedData_15(lis_io_sortedData_15),
    .io_sortedData_16(lis_io_sortedData_16),
    .io_sortedData_17(lis_io_sortedData_17),
    .io_sortedData_18(lis_io_sortedData_18),
    .io_sortedData_19(lis_io_sortedData_19),
    .io_sortedData_20(lis_io_sortedData_20),
    .io_sortedData_21(lis_io_sortedData_21),
    .io_sortedData_22(lis_io_sortedData_22),
    .io_sortedData_23(lis_io_sortedData_23),
    .io_sorterFull(lis_io_sorterFull),
    .io_sorterEmpty(lis_io_sorterEmpty),
    .io_lisSize(lis_io_lisSize),
    .io_discardPos(lis_io_discardPos)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_stream_in_bits_data; // @[LISDspBlock.scala 71:44]
  assign _GEN_0 = lis_io_sortedData_0; // @[LISDspBlock.scala 92:82]
  assign _GEN_1 = 5'h1 == sendOnOutput ? $signed(lis_io_sortedData_1) : $signed(_GEN_0); // @[LISDspBlock.scala 92:82]
  assign _GEN_2 = 5'h2 == sendOnOutput ? $signed(lis_io_sortedData_2) : $signed(_GEN_1); // @[LISDspBlock.scala 92:82]
  assign _GEN_3 = 5'h3 == sendOnOutput ? $signed(lis_io_sortedData_3) : $signed(_GEN_2); // @[LISDspBlock.scala 92:82]
  assign _GEN_4 = 5'h4 == sendOnOutput ? $signed(lis_io_sortedData_4) : $signed(_GEN_3); // @[LISDspBlock.scala 92:82]
  assign _GEN_5 = 5'h5 == sendOnOutput ? $signed(lis_io_sortedData_5) : $signed(_GEN_4); // @[LISDspBlock.scala 92:82]
  assign _GEN_6 = 5'h6 == sendOnOutput ? $signed(lis_io_sortedData_6) : $signed(_GEN_5); // @[LISDspBlock.scala 92:82]
  assign _GEN_7 = 5'h7 == sendOnOutput ? $signed(lis_io_sortedData_7) : $signed(_GEN_6); // @[LISDspBlock.scala 92:82]
  assign _GEN_8 = 5'h8 == sendOnOutput ? $signed(lis_io_sortedData_8) : $signed(_GEN_7); // @[LISDspBlock.scala 92:82]
  assign _GEN_9 = 5'h9 == sendOnOutput ? $signed(lis_io_sortedData_9) : $signed(_GEN_8); // @[LISDspBlock.scala 92:82]
  assign _GEN_10 = 5'ha == sendOnOutput ? $signed(lis_io_sortedData_10) : $signed(_GEN_9); // @[LISDspBlock.scala 92:82]
  assign _GEN_11 = 5'hb == sendOnOutput ? $signed(lis_io_sortedData_11) : $signed(_GEN_10); // @[LISDspBlock.scala 92:82]
  assign _GEN_12 = 5'hc == sendOnOutput ? $signed(lis_io_sortedData_12) : $signed(_GEN_11); // @[LISDspBlock.scala 92:82]
  assign _GEN_13 = 5'hd == sendOnOutput ? $signed(lis_io_sortedData_13) : $signed(_GEN_12); // @[LISDspBlock.scala 92:82]
  assign _GEN_14 = 5'he == sendOnOutput ? $signed(lis_io_sortedData_14) : $signed(_GEN_13); // @[LISDspBlock.scala 92:82]
  assign _GEN_15 = 5'hf == sendOnOutput ? $signed(lis_io_sortedData_15) : $signed(_GEN_14); // @[LISDspBlock.scala 92:82]
  assign _GEN_16 = 5'h10 == sendOnOutput ? $signed(lis_io_sortedData_16) : $signed(_GEN_15); // @[LISDspBlock.scala 92:82]
  assign _GEN_17 = 5'h11 == sendOnOutput ? $signed(lis_io_sortedData_17) : $signed(_GEN_16); // @[LISDspBlock.scala 92:82]
  assign _GEN_18 = 5'h12 == sendOnOutput ? $signed(lis_io_sortedData_18) : $signed(_GEN_17); // @[LISDspBlock.scala 92:82]
  assign _GEN_19 = 5'h13 == sendOnOutput ? $signed(lis_io_sortedData_19) : $signed(_GEN_18); // @[LISDspBlock.scala 92:82]
  assign _GEN_20 = 5'h14 == sendOnOutput ? $signed(lis_io_sortedData_20) : $signed(_GEN_19); // @[LISDspBlock.scala 92:82]
  assign _GEN_21 = 5'h15 == sendOnOutput ? $signed(lis_io_sortedData_21) : $signed(_GEN_20); // @[LISDspBlock.scala 92:82]
  assign _GEN_22 = 5'h16 == sendOnOutput ? $signed(lis_io_sortedData_22) : $signed(_GEN_21); // @[LISDspBlock.scala 92:82]
  assign _T_4 = 5'h17 == sendOnOutput ? $signed(lis_io_sortedData_23) : $signed(_GEN_22); // @[LISDspBlock.scala 92:82]
  assign _T_7 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_8 = auto_mem_in_ar_valid | _T_7; // @[RegisterRouter.scala 40:26]
  assign _T_9 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_52_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_16 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_281 = {_T_16[4],_T_16[3],_T_16[2]}; // @[Cat.scala 29:58]
  assign _T_56 = _T_16[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_64 = _T_56 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_10 = _T_52_ready & _T_9; // @[RegisterRouter.scala 42:26]
  assign _T_19 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_21 = _T_19 | 2'h1; // @[Misc.scala 200:81]
  assign _T_22 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_25 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_27 = _T_21[1] & _T_25; // @[Misc.scala 213:38]
  assign _T_28 = _T_22 | _T_27; // @[Misc.scala 213:29]
  assign _T_30 = _T_21[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_31 = _T_22 | _T_30; // @[Misc.scala 213:29]
  assign _T_34 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_35 = _T_25 & _T_34; // @[Misc.scala 212:27]
  assign _T_36 = _T_21[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = _T_25 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_39 = _T_21[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & _T_34; // @[Misc.scala 212:27]
  assign _T_42 = _T_21[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_31 | _T_42; // @[Misc.scala 213:29]
  assign _T_44 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_45 = _T_21[0] & _T_44; // @[Misc.scala 213:38]
  assign _T_46 = _T_31 | _T_45; // @[Misc.scala 213:29]
  assign _T_49 = {_T_46,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  assign _T_51 = auto_mem_in_ar_valid ? _T_49 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_51[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_51[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_51[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_51[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_300 = _T_8 & _T_52_ready; // @[RegisterRouter.scala 59:16]
  assign _T_282 = 8'h1 << _T_281; // @[OneHot.scala 58:35]
  assign _T_347 = _T_300 & _T_9; // @[RegisterRouter.scala 59:16]
  assign _T_349 = _T_347 & _T_282[0]; // @[RegisterRouter.scala 59:16]
  assign _T_350 = _T_349 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_350 & _T_89[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_24 = _T_115 ? auto_mem_in_w_bits_data[0] : sortDir; // @[RegField.scala 134:88]
  assign _T_154 = _T_89[4:0] == 5'h1f; // @[RegisterRouter.scala 59:16]
  assign _T_354 = _T_347 & _T_282[1]; // @[RegisterRouter.scala 59:16]
  assign _T_355 = _T_354 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_355 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _T_359 = _T_347 & _T_282[2]; // @[RegisterRouter.scala 59:16]
  assign _T_360 = _T_359 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_207 = _T_360 & _T_89[0]; // @[RegisterRouter.scala 59:16]
  assign _T_364 = _T_347 & _T_282[3]; // @[RegisterRouter.scala 59:16]
  assign _T_365 = _T_364 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_230 = _T_365 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _T_369 = _T_347 & _T_282[4]; // @[RegisterRouter.scala 59:16]
  assign _T_370 = _T_369 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_253 = _T_370 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _GEN_62 = 3'h1 == _T_281 ? _T_64 : _T_64; // @[MuxLiteral.scala 48:10]
  assign _GEN_63 = 3'h2 == _T_281 ? _T_64 : _GEN_62; // @[MuxLiteral.scala 48:10]
  assign _GEN_64 = 3'h3 == _T_281 ? _T_64 : _GEN_63; // @[MuxLiteral.scala 48:10]
  assign _GEN_65 = 3'h4 == _T_281 ? _T_64 : _GEN_64; // @[MuxLiteral.scala 48:10]
  assign _GEN_66 = 3'h5 == _T_281 ? _T_64 : _GEN_65; // @[MuxLiteral.scala 48:10]
  assign _GEN_67 = 3'h6 == _T_281 ? _T_64 : _GEN_66; // @[MuxLiteral.scala 48:10]
  assign _GEN_77 = 3'h7 == _T_281; // @[MuxLiteral.scala 48:10]
  assign _GEN_68 = _GEN_77 | _GEN_67; // @[MuxLiteral.scala 48:10]
  assign _T_492_0 = {{4'd0}, sortDir}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_70 = 3'h1 == _T_281 ? lisSize : _T_492_0; // @[MuxLiteral.scala 48:10]
  assign _T_492_2 = {{4'd0}, flushData}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_71 = 3'h2 == _T_281 ? _T_492_2 : _GEN_70; // @[MuxLiteral.scala 48:10]
  assign _GEN_72 = 3'h3 == _T_281 ? discardPos : _GEN_71; // @[MuxLiteral.scala 48:10]
  assign _GEN_73 = 3'h4 == _T_281 ? sendOnOutput : _GEN_72; // @[MuxLiteral.scala 48:10]
  assign _T_492_5 = {{4'd0}, sorterFull}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_74 = 3'h5 == _T_281 ? _T_492_5 : _GEN_73; // @[MuxLiteral.scala 48:10]
  assign _T_492_6 = {{4'd0}, sorterEmpty}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_75 = 3'h6 == _T_281 ? _T_492_6 : _GEN_74; // @[MuxLiteral.scala 48:10]
  assign _GEN_76 = 3'h7 == _T_281 ? 5'h0 : _GEN_75; // @[MuxLiteral.scala 48:10]
  assign _T_494 = _GEN_68 ? _GEN_76 : 5'h0; // @[RegisterRouter.scala 59:16]
  assign _T_495_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_495_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_498 = ~_T_495_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_10 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_10 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_495_valid & _T_498; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_495_valid & _T_495_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = lis_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = lis_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {lis_io_out_bits,_T_4}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = lis_io_lastOut; // @[LazyModule.scala 173:49]
  assign lis_clock = clock;
  assign lis_reset = reset;
  assign lis_io_in_valid = auto_stream_in_valid; // @[LISDspBlock.scala 70:21]
  assign lis_io_in_bits = _T_2[15:0]; // @[LISDspBlock.scala 71:20]
  assign lis_io_lastIn = auto_stream_in_bits_last; // @[LISDspBlock.scala 69:19]
  assign lis_io_out_ready = auto_stream_out_ready; // @[LISDspBlock.scala 91:22]
  assign lis_io_lisSize = {{1'd0}, lisSize}; // @[LISDspBlock.scala 79:26]
  assign lis_io_discardPos = discardPos; // @[LISDspBlock.scala 85:29]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_7; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{27'd0}, _T_494}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_495_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sortDir = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flushData = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  discardPos = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sendOnOutput = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  lisSize = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sorterFull = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sorterEmpty = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sortDir <= reset | _GEN_24;
    if (reset) begin
      flushData <= 1'h0;
    end else if (_T_207) begin
      flushData <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      discardPos <= 5'h0;
    end else if (_T_230) begin
      discardPos <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      sendOnOutput <= 5'h0;
    end else if (_T_253) begin
      sendOnOutput <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      lisSize <= 5'h18;
    end else if (_T_161) begin
      lisSize <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      sorterFull <= 1'h0;
    end else begin
      sorterFull <= lis_io_sorterFull;
    end
    sorterEmpty <= reset | lis_io_sorterEmpty;
  end
endmodule
module LinearSorter_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [15:0] io_in_bits,
  input         io_lastIn,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits,
  output        io_lastOut,
  output [15:0] io_sortedData_0,
  output [15:0] io_sortedData_1,
  output [15:0] io_sortedData_2,
  output [15:0] io_sortedData_3,
  output [15:0] io_sortedData_4,
  output [15:0] io_sortedData_5,
  output [15:0] io_sortedData_6,
  output [15:0] io_sortedData_7,
  output [15:0] io_sortedData_8,
  output [15:0] io_sortedData_9,
  output [15:0] io_sortedData_10,
  output [15:0] io_sortedData_11,
  output [15:0] io_sortedData_12,
  output [15:0] io_sortedData_13,
  output [15:0] io_sortedData_14,
  output [15:0] io_sortedData_15,
  output [15:0] io_sortedData_16,
  output [15:0] io_sortedData_17,
  output [15:0] io_sortedData_18,
  output [15:0] io_sortedData_19,
  output [15:0] io_sortedData_20,
  output [15:0] io_sortedData_21,
  output [15:0] io_sortedData_22,
  output [15:0] io_sortedData_23,
  output        io_sorterFull,
  output        io_sorterEmpty,
  input  [5:0]  io_lisSize
);
  wire  PEChain_0_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_0_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_0_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_0_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_1_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_1_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_1_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_2_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_2_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_2_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_3_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_3_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_3_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_4_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_4_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_4_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_5_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_5_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_5_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_6_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_6_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_6_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_7_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_7_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_7_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_8_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_8_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_8_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_9_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_9_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_9_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_10_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_10_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_10_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_11_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_11_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_11_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_12_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_12_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_12_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_13_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_13_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_13_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_14_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_14_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_14_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_15_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_15_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_15_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_16_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_16_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_16_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_17_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_17_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_17_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_18_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_18_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_18_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_19_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_19_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_19_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_20_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_20_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_20_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_21_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_21_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_21_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_22_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_rightNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_rightNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_inData; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_rightPropDiscard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_22_io_rightOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_22_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_clock; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_reset; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_enableSort; // @[LinearSorter.scala 143:24]
  wire [1:0] PEChain_23_io_state; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_leftNBR_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_leftNBR_compRes; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_currCell_data; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_currCell_compRes; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_lastCell; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_active; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_discard; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_inData; // @[LinearSorter.scala 143:24]
  wire [15:0] PEChain_23_io_leftOutData; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_currDiscard; // @[LinearSorter.scala 143:24]
  wire  PEChain_23_io_toLeftPropDiscard; // @[LinearSorter.scala 143:24]
  reg  initialInDone; // @[LinearSorter.scala 67:30]
  reg [31:0] _RAND_0;
  reg [4:0] cntInData; // @[LinearSorter.scala 68:26]
  reg [31:0] _RAND_1;
  reg [1:0] state; // @[LinearSorter.scala 78:22]
  reg [31:0] _RAND_2;
  reg [5:0] lisSizeReg; // @[LinearSorter.scala 81:27]
  reg [31:0] _RAND_3;
  wire [5:0] _T_1; // @[LinearSorter.scala 86:43]
  wire  _T_96; // @[Decoupled.scala 40:37]
  wire [4:0] _T_98; // @[LinearSorter.scala 92:28]
  wire  _T_99; // @[LinearSorter.scala 94:20]
  wire [5:0] _GEN_111; // @[LinearSorter.scala 98:19]
  wire  _T_102; // @[LinearSorter.scala 98:19]
  wire  _T_104; // @[LinearSorter.scala 98:42]
  wire  _T_113; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_7; // @[LinearSorter.scala 117:27]
  wire  _T_115; // @[Conditional.scala 37:30]
  wire  fireLastIn; // @[LinearSorter.scala 111:30]
  wire [1:0] _GEN_8; // @[LinearSorter.scala 120:62]
  wire  _T_117; // @[Conditional.scala 37:30]
  reg [4:0] cntOutData; // @[LISutil.scala 10:33]
  reg [31:0] _RAND_4;
  wire [5:0] _GEN_112; // @[LinearSorter.scala 125:28]
  wire  _T_120; // @[LinearSorter.scala 125:28]
  wire [1:0] _GEN_9; // @[LinearSorter.scala 125:50]
  wire [1:0] _GEN_10; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_11; // @[Conditional.scala 39:67]
  wire [1:0] state_next; // @[Conditional.scala 40:58]
  wire  _T_105; // @[LinearSorter.scala 101:25]
  wire  _GEN_2; // @[LinearSorter.scala 101:36]
  wire  _GEN_3; // @[LinearSorter.scala 98:59]
  wire  _T_106; // @[LinearSorter.scala 106:29]
  wire  _T_107; // @[LinearSorter.scala 106:54]
  wire  enable; // @[LinearSorter.scala 106:45]
  wire  _T_109; // @[LISutil.scala 13:24]
  wire [4:0] _T_111; // @[LISutil.scala 14:22]
  wire  _T_121; // @[LinearSorter.scala 137:33]
  wire [15:0] outputData_0; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] outputData_1; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_16; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_2; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_17; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_3; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_18; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_4; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_19; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_5; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_20; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_6; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_21; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_7; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_22; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_8; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_23; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_9; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_24; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_10; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_25; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_11; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_26; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_12; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_27; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_13; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_28; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_14; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_29; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_15; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_30; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_16; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_31; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_17; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_32; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_18; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_33; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_19; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_34; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_20; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_35; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_21; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_36; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_22; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_37; // @[LinearSorter.scala 137:21]
  wire [15:0] outputData_23; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  wire [15:0] _GEN_38; // @[LinearSorter.scala 137:21]
  wire  _T_136; // @[LinearSorter.scala 168:63]
  wire  discardSignals_2; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_1; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_0; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_5; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_4; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_3; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [5:0] _T_372; // @[LinearSorter.scala 177:50]
  wire  discardSignals_8; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_7; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_6; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_11; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_10; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_9; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [11:0] _T_378; // @[LinearSorter.scala 177:50]
  wire  discardSignals_14; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_13; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_12; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_17; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_16; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_15; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [5:0] _T_383; // @[LinearSorter.scala 177:50]
  wire  discardSignals_20; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_19; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_18; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_23; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_22; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire  discardSignals_21; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  wire [23:0] _T_390; // @[LinearSorter.scala 177:50]
  wire [4:0] _T_415; // @[Mux.scala 47:69]
  wire [4:0] _T_416; // @[Mux.scala 47:69]
  wire [4:0] _T_417; // @[Mux.scala 47:69]
  wire [4:0] _T_418; // @[Mux.scala 47:69]
  wire [4:0] _T_419; // @[Mux.scala 47:69]
  wire [4:0] _T_420; // @[Mux.scala 47:69]
  wire [4:0] _T_421; // @[Mux.scala 47:69]
  wire [4:0] _T_422; // @[Mux.scala 47:69]
  wire [4:0] _T_423; // @[Mux.scala 47:69]
  wire [4:0] _T_424; // @[Mux.scala 47:69]
  wire [4:0] _T_425; // @[Mux.scala 47:69]
  wire [4:0] _T_426; // @[Mux.scala 47:69]
  wire [4:0] _T_427; // @[Mux.scala 47:69]
  wire [4:0] _T_428; // @[Mux.scala 47:69]
  wire [4:0] _T_429; // @[Mux.scala 47:69]
  wire [4:0] _T_430; // @[Mux.scala 47:69]
  wire [4:0] _T_431; // @[Mux.scala 47:69]
  wire [4:0] _T_432; // @[Mux.scala 47:69]
  wire [4:0] _T_433; // @[Mux.scala 47:69]
  wire [4:0] _T_434; // @[Mux.scala 47:69]
  wire [4:0] _T_435; // @[Mux.scala 47:69]
  wire [4:0] _T_436; // @[Mux.scala 47:69]
  wire [4:0] getDiscarded; // @[Mux.scala 47:69]
  wire  _T_438; // @[LinearSorter.scala 199:49]
  wire [15:0] _GEN_88; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_89; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_90; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_91; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_92; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_93; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_94; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_95; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_96; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_97; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_98; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_99; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_100; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_101; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_102; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_103; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_104; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_105; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_106; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_107; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_108; // @[LinearSorter.scala 206:15]
  wire [15:0] _GEN_109; // @[LinearSorter.scala 206:15]
  wire  _T_444; // @[LinearSorter.scala 208:18]
  wire  _T_446; // @[LinearSorter.scala 208:49]
  wire  _T_448; // @[LinearSorter.scala 209:33]
  PE_24 PEChain_0 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_0_clock),
    .reset(PEChain_0_reset),
    .io_enableSort(PEChain_0_io_enableSort),
    .io_state(PEChain_0_io_state),
    .io_rightNBR_data(PEChain_0_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_0_io_rightNBR_compRes),
    .io_currCell_data(PEChain_0_io_currCell_data),
    .io_currCell_compRes(PEChain_0_io_currCell_compRes),
    .io_lastCell(PEChain_0_io_lastCell),
    .io_discard(PEChain_0_io_discard),
    .io_inData(PEChain_0_io_inData),
    .io_rightPropDiscard(PEChain_0_io_rightPropDiscard),
    .io_rightOutData(PEChain_0_io_rightOutData),
    .io_currDiscard(PEChain_0_io_currDiscard)
  );
  PE_25 PEChain_1 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_1_clock),
    .reset(PEChain_1_reset),
    .io_enableSort(PEChain_1_io_enableSort),
    .io_state(PEChain_1_io_state),
    .io_leftNBR_data(PEChain_1_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_1_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_1_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_1_io_rightNBR_compRes),
    .io_currCell_data(PEChain_1_io_currCell_data),
    .io_currCell_compRes(PEChain_1_io_currCell_compRes),
    .io_lastCell(PEChain_1_io_lastCell),
    .io_active(PEChain_1_io_active),
    .io_discard(PEChain_1_io_discard),
    .io_inData(PEChain_1_io_inData),
    .io_rightPropDiscard(PEChain_1_io_rightPropDiscard),
    .io_leftOutData(PEChain_1_io_leftOutData),
    .io_rightOutData(PEChain_1_io_rightOutData),
    .io_currDiscard(PEChain_1_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_1_io_toLeftPropDiscard)
  );
  PE_26 PEChain_2 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_2_clock),
    .reset(PEChain_2_reset),
    .io_enableSort(PEChain_2_io_enableSort),
    .io_state(PEChain_2_io_state),
    .io_leftNBR_data(PEChain_2_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_2_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_2_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_2_io_rightNBR_compRes),
    .io_currCell_data(PEChain_2_io_currCell_data),
    .io_currCell_compRes(PEChain_2_io_currCell_compRes),
    .io_lastCell(PEChain_2_io_lastCell),
    .io_active(PEChain_2_io_active),
    .io_discard(PEChain_2_io_discard),
    .io_inData(PEChain_2_io_inData),
    .io_rightPropDiscard(PEChain_2_io_rightPropDiscard),
    .io_leftOutData(PEChain_2_io_leftOutData),
    .io_rightOutData(PEChain_2_io_rightOutData),
    .io_currDiscard(PEChain_2_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_2_io_toLeftPropDiscard)
  );
  PE_27 PEChain_3 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_3_clock),
    .reset(PEChain_3_reset),
    .io_enableSort(PEChain_3_io_enableSort),
    .io_state(PEChain_3_io_state),
    .io_leftNBR_data(PEChain_3_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_3_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_3_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_3_io_rightNBR_compRes),
    .io_currCell_data(PEChain_3_io_currCell_data),
    .io_currCell_compRes(PEChain_3_io_currCell_compRes),
    .io_lastCell(PEChain_3_io_lastCell),
    .io_active(PEChain_3_io_active),
    .io_discard(PEChain_3_io_discard),
    .io_inData(PEChain_3_io_inData),
    .io_rightPropDiscard(PEChain_3_io_rightPropDiscard),
    .io_leftOutData(PEChain_3_io_leftOutData),
    .io_rightOutData(PEChain_3_io_rightOutData),
    .io_currDiscard(PEChain_3_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_3_io_toLeftPropDiscard)
  );
  PE_28 PEChain_4 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_4_clock),
    .reset(PEChain_4_reset),
    .io_enableSort(PEChain_4_io_enableSort),
    .io_state(PEChain_4_io_state),
    .io_leftNBR_data(PEChain_4_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_4_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_4_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_4_io_rightNBR_compRes),
    .io_currCell_data(PEChain_4_io_currCell_data),
    .io_currCell_compRes(PEChain_4_io_currCell_compRes),
    .io_lastCell(PEChain_4_io_lastCell),
    .io_active(PEChain_4_io_active),
    .io_discard(PEChain_4_io_discard),
    .io_inData(PEChain_4_io_inData),
    .io_rightPropDiscard(PEChain_4_io_rightPropDiscard),
    .io_leftOutData(PEChain_4_io_leftOutData),
    .io_rightOutData(PEChain_4_io_rightOutData),
    .io_currDiscard(PEChain_4_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_4_io_toLeftPropDiscard)
  );
  PE_29 PEChain_5 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_5_clock),
    .reset(PEChain_5_reset),
    .io_enableSort(PEChain_5_io_enableSort),
    .io_state(PEChain_5_io_state),
    .io_leftNBR_data(PEChain_5_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_5_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_5_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_5_io_rightNBR_compRes),
    .io_currCell_data(PEChain_5_io_currCell_data),
    .io_currCell_compRes(PEChain_5_io_currCell_compRes),
    .io_lastCell(PEChain_5_io_lastCell),
    .io_active(PEChain_5_io_active),
    .io_discard(PEChain_5_io_discard),
    .io_inData(PEChain_5_io_inData),
    .io_rightPropDiscard(PEChain_5_io_rightPropDiscard),
    .io_leftOutData(PEChain_5_io_leftOutData),
    .io_rightOutData(PEChain_5_io_rightOutData),
    .io_currDiscard(PEChain_5_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_5_io_toLeftPropDiscard)
  );
  PE_30 PEChain_6 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_6_clock),
    .reset(PEChain_6_reset),
    .io_enableSort(PEChain_6_io_enableSort),
    .io_state(PEChain_6_io_state),
    .io_leftNBR_data(PEChain_6_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_6_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_6_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_6_io_rightNBR_compRes),
    .io_currCell_data(PEChain_6_io_currCell_data),
    .io_currCell_compRes(PEChain_6_io_currCell_compRes),
    .io_lastCell(PEChain_6_io_lastCell),
    .io_active(PEChain_6_io_active),
    .io_discard(PEChain_6_io_discard),
    .io_inData(PEChain_6_io_inData),
    .io_rightPropDiscard(PEChain_6_io_rightPropDiscard),
    .io_leftOutData(PEChain_6_io_leftOutData),
    .io_rightOutData(PEChain_6_io_rightOutData),
    .io_currDiscard(PEChain_6_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_6_io_toLeftPropDiscard)
  );
  PE_31 PEChain_7 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_7_clock),
    .reset(PEChain_7_reset),
    .io_enableSort(PEChain_7_io_enableSort),
    .io_state(PEChain_7_io_state),
    .io_leftNBR_data(PEChain_7_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_7_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_7_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_7_io_rightNBR_compRes),
    .io_currCell_data(PEChain_7_io_currCell_data),
    .io_currCell_compRes(PEChain_7_io_currCell_compRes),
    .io_lastCell(PEChain_7_io_lastCell),
    .io_active(PEChain_7_io_active),
    .io_discard(PEChain_7_io_discard),
    .io_inData(PEChain_7_io_inData),
    .io_rightPropDiscard(PEChain_7_io_rightPropDiscard),
    .io_leftOutData(PEChain_7_io_leftOutData),
    .io_rightOutData(PEChain_7_io_rightOutData),
    .io_currDiscard(PEChain_7_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_7_io_toLeftPropDiscard)
  );
  PE_32 PEChain_8 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_8_clock),
    .reset(PEChain_8_reset),
    .io_enableSort(PEChain_8_io_enableSort),
    .io_state(PEChain_8_io_state),
    .io_leftNBR_data(PEChain_8_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_8_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_8_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_8_io_rightNBR_compRes),
    .io_currCell_data(PEChain_8_io_currCell_data),
    .io_currCell_compRes(PEChain_8_io_currCell_compRes),
    .io_lastCell(PEChain_8_io_lastCell),
    .io_active(PEChain_8_io_active),
    .io_discard(PEChain_8_io_discard),
    .io_inData(PEChain_8_io_inData),
    .io_rightPropDiscard(PEChain_8_io_rightPropDiscard),
    .io_leftOutData(PEChain_8_io_leftOutData),
    .io_rightOutData(PEChain_8_io_rightOutData),
    .io_currDiscard(PEChain_8_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_8_io_toLeftPropDiscard)
  );
  PE_33 PEChain_9 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_9_clock),
    .reset(PEChain_9_reset),
    .io_enableSort(PEChain_9_io_enableSort),
    .io_state(PEChain_9_io_state),
    .io_leftNBR_data(PEChain_9_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_9_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_9_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_9_io_rightNBR_compRes),
    .io_currCell_data(PEChain_9_io_currCell_data),
    .io_currCell_compRes(PEChain_9_io_currCell_compRes),
    .io_lastCell(PEChain_9_io_lastCell),
    .io_active(PEChain_9_io_active),
    .io_discard(PEChain_9_io_discard),
    .io_inData(PEChain_9_io_inData),
    .io_rightPropDiscard(PEChain_9_io_rightPropDiscard),
    .io_leftOutData(PEChain_9_io_leftOutData),
    .io_rightOutData(PEChain_9_io_rightOutData),
    .io_currDiscard(PEChain_9_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_9_io_toLeftPropDiscard)
  );
  PE_34 PEChain_10 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_10_clock),
    .reset(PEChain_10_reset),
    .io_enableSort(PEChain_10_io_enableSort),
    .io_state(PEChain_10_io_state),
    .io_leftNBR_data(PEChain_10_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_10_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_10_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_10_io_rightNBR_compRes),
    .io_currCell_data(PEChain_10_io_currCell_data),
    .io_currCell_compRes(PEChain_10_io_currCell_compRes),
    .io_lastCell(PEChain_10_io_lastCell),
    .io_active(PEChain_10_io_active),
    .io_discard(PEChain_10_io_discard),
    .io_inData(PEChain_10_io_inData),
    .io_rightPropDiscard(PEChain_10_io_rightPropDiscard),
    .io_leftOutData(PEChain_10_io_leftOutData),
    .io_rightOutData(PEChain_10_io_rightOutData),
    .io_currDiscard(PEChain_10_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_10_io_toLeftPropDiscard)
  );
  PE_35 PEChain_11 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_11_clock),
    .reset(PEChain_11_reset),
    .io_enableSort(PEChain_11_io_enableSort),
    .io_state(PEChain_11_io_state),
    .io_leftNBR_data(PEChain_11_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_11_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_11_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_11_io_rightNBR_compRes),
    .io_currCell_data(PEChain_11_io_currCell_data),
    .io_currCell_compRes(PEChain_11_io_currCell_compRes),
    .io_lastCell(PEChain_11_io_lastCell),
    .io_active(PEChain_11_io_active),
    .io_discard(PEChain_11_io_discard),
    .io_inData(PEChain_11_io_inData),
    .io_rightPropDiscard(PEChain_11_io_rightPropDiscard),
    .io_leftOutData(PEChain_11_io_leftOutData),
    .io_rightOutData(PEChain_11_io_rightOutData),
    .io_currDiscard(PEChain_11_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_11_io_toLeftPropDiscard)
  );
  PE_36 PEChain_12 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_12_clock),
    .reset(PEChain_12_reset),
    .io_enableSort(PEChain_12_io_enableSort),
    .io_state(PEChain_12_io_state),
    .io_leftNBR_data(PEChain_12_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_12_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_12_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_12_io_rightNBR_compRes),
    .io_currCell_data(PEChain_12_io_currCell_data),
    .io_currCell_compRes(PEChain_12_io_currCell_compRes),
    .io_lastCell(PEChain_12_io_lastCell),
    .io_active(PEChain_12_io_active),
    .io_discard(PEChain_12_io_discard),
    .io_inData(PEChain_12_io_inData),
    .io_rightPropDiscard(PEChain_12_io_rightPropDiscard),
    .io_leftOutData(PEChain_12_io_leftOutData),
    .io_rightOutData(PEChain_12_io_rightOutData),
    .io_currDiscard(PEChain_12_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_12_io_toLeftPropDiscard)
  );
  PE_37 PEChain_13 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_13_clock),
    .reset(PEChain_13_reset),
    .io_enableSort(PEChain_13_io_enableSort),
    .io_state(PEChain_13_io_state),
    .io_leftNBR_data(PEChain_13_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_13_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_13_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_13_io_rightNBR_compRes),
    .io_currCell_data(PEChain_13_io_currCell_data),
    .io_currCell_compRes(PEChain_13_io_currCell_compRes),
    .io_lastCell(PEChain_13_io_lastCell),
    .io_active(PEChain_13_io_active),
    .io_discard(PEChain_13_io_discard),
    .io_inData(PEChain_13_io_inData),
    .io_rightPropDiscard(PEChain_13_io_rightPropDiscard),
    .io_leftOutData(PEChain_13_io_leftOutData),
    .io_rightOutData(PEChain_13_io_rightOutData),
    .io_currDiscard(PEChain_13_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_13_io_toLeftPropDiscard)
  );
  PE_38 PEChain_14 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_14_clock),
    .reset(PEChain_14_reset),
    .io_enableSort(PEChain_14_io_enableSort),
    .io_state(PEChain_14_io_state),
    .io_leftNBR_data(PEChain_14_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_14_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_14_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_14_io_rightNBR_compRes),
    .io_currCell_data(PEChain_14_io_currCell_data),
    .io_currCell_compRes(PEChain_14_io_currCell_compRes),
    .io_lastCell(PEChain_14_io_lastCell),
    .io_active(PEChain_14_io_active),
    .io_discard(PEChain_14_io_discard),
    .io_inData(PEChain_14_io_inData),
    .io_rightPropDiscard(PEChain_14_io_rightPropDiscard),
    .io_leftOutData(PEChain_14_io_leftOutData),
    .io_rightOutData(PEChain_14_io_rightOutData),
    .io_currDiscard(PEChain_14_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_14_io_toLeftPropDiscard)
  );
  PE_39 PEChain_15 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_15_clock),
    .reset(PEChain_15_reset),
    .io_enableSort(PEChain_15_io_enableSort),
    .io_state(PEChain_15_io_state),
    .io_leftNBR_data(PEChain_15_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_15_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_15_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_15_io_rightNBR_compRes),
    .io_currCell_data(PEChain_15_io_currCell_data),
    .io_currCell_compRes(PEChain_15_io_currCell_compRes),
    .io_lastCell(PEChain_15_io_lastCell),
    .io_active(PEChain_15_io_active),
    .io_discard(PEChain_15_io_discard),
    .io_inData(PEChain_15_io_inData),
    .io_rightPropDiscard(PEChain_15_io_rightPropDiscard),
    .io_leftOutData(PEChain_15_io_leftOutData),
    .io_rightOutData(PEChain_15_io_rightOutData),
    .io_currDiscard(PEChain_15_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_15_io_toLeftPropDiscard)
  );
  PE_40 PEChain_16 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_16_clock),
    .reset(PEChain_16_reset),
    .io_enableSort(PEChain_16_io_enableSort),
    .io_state(PEChain_16_io_state),
    .io_leftNBR_data(PEChain_16_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_16_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_16_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_16_io_rightNBR_compRes),
    .io_currCell_data(PEChain_16_io_currCell_data),
    .io_currCell_compRes(PEChain_16_io_currCell_compRes),
    .io_lastCell(PEChain_16_io_lastCell),
    .io_active(PEChain_16_io_active),
    .io_discard(PEChain_16_io_discard),
    .io_inData(PEChain_16_io_inData),
    .io_rightPropDiscard(PEChain_16_io_rightPropDiscard),
    .io_leftOutData(PEChain_16_io_leftOutData),
    .io_rightOutData(PEChain_16_io_rightOutData),
    .io_currDiscard(PEChain_16_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_16_io_toLeftPropDiscard)
  );
  PE_41 PEChain_17 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_17_clock),
    .reset(PEChain_17_reset),
    .io_enableSort(PEChain_17_io_enableSort),
    .io_state(PEChain_17_io_state),
    .io_leftNBR_data(PEChain_17_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_17_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_17_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_17_io_rightNBR_compRes),
    .io_currCell_data(PEChain_17_io_currCell_data),
    .io_currCell_compRes(PEChain_17_io_currCell_compRes),
    .io_lastCell(PEChain_17_io_lastCell),
    .io_active(PEChain_17_io_active),
    .io_discard(PEChain_17_io_discard),
    .io_inData(PEChain_17_io_inData),
    .io_rightPropDiscard(PEChain_17_io_rightPropDiscard),
    .io_leftOutData(PEChain_17_io_leftOutData),
    .io_rightOutData(PEChain_17_io_rightOutData),
    .io_currDiscard(PEChain_17_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_17_io_toLeftPropDiscard)
  );
  PE_42 PEChain_18 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_18_clock),
    .reset(PEChain_18_reset),
    .io_enableSort(PEChain_18_io_enableSort),
    .io_state(PEChain_18_io_state),
    .io_leftNBR_data(PEChain_18_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_18_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_18_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_18_io_rightNBR_compRes),
    .io_currCell_data(PEChain_18_io_currCell_data),
    .io_currCell_compRes(PEChain_18_io_currCell_compRes),
    .io_lastCell(PEChain_18_io_lastCell),
    .io_active(PEChain_18_io_active),
    .io_discard(PEChain_18_io_discard),
    .io_inData(PEChain_18_io_inData),
    .io_rightPropDiscard(PEChain_18_io_rightPropDiscard),
    .io_leftOutData(PEChain_18_io_leftOutData),
    .io_rightOutData(PEChain_18_io_rightOutData),
    .io_currDiscard(PEChain_18_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_18_io_toLeftPropDiscard)
  );
  PE_43 PEChain_19 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_19_clock),
    .reset(PEChain_19_reset),
    .io_enableSort(PEChain_19_io_enableSort),
    .io_state(PEChain_19_io_state),
    .io_leftNBR_data(PEChain_19_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_19_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_19_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_19_io_rightNBR_compRes),
    .io_currCell_data(PEChain_19_io_currCell_data),
    .io_currCell_compRes(PEChain_19_io_currCell_compRes),
    .io_lastCell(PEChain_19_io_lastCell),
    .io_active(PEChain_19_io_active),
    .io_discard(PEChain_19_io_discard),
    .io_inData(PEChain_19_io_inData),
    .io_rightPropDiscard(PEChain_19_io_rightPropDiscard),
    .io_leftOutData(PEChain_19_io_leftOutData),
    .io_rightOutData(PEChain_19_io_rightOutData),
    .io_currDiscard(PEChain_19_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_19_io_toLeftPropDiscard)
  );
  PE_44 PEChain_20 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_20_clock),
    .reset(PEChain_20_reset),
    .io_enableSort(PEChain_20_io_enableSort),
    .io_state(PEChain_20_io_state),
    .io_leftNBR_data(PEChain_20_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_20_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_20_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_20_io_rightNBR_compRes),
    .io_currCell_data(PEChain_20_io_currCell_data),
    .io_currCell_compRes(PEChain_20_io_currCell_compRes),
    .io_lastCell(PEChain_20_io_lastCell),
    .io_active(PEChain_20_io_active),
    .io_discard(PEChain_20_io_discard),
    .io_inData(PEChain_20_io_inData),
    .io_rightPropDiscard(PEChain_20_io_rightPropDiscard),
    .io_leftOutData(PEChain_20_io_leftOutData),
    .io_rightOutData(PEChain_20_io_rightOutData),
    .io_currDiscard(PEChain_20_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_20_io_toLeftPropDiscard)
  );
  PE_45 PEChain_21 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_21_clock),
    .reset(PEChain_21_reset),
    .io_enableSort(PEChain_21_io_enableSort),
    .io_state(PEChain_21_io_state),
    .io_leftNBR_data(PEChain_21_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_21_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_21_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_21_io_rightNBR_compRes),
    .io_currCell_data(PEChain_21_io_currCell_data),
    .io_currCell_compRes(PEChain_21_io_currCell_compRes),
    .io_lastCell(PEChain_21_io_lastCell),
    .io_active(PEChain_21_io_active),
    .io_discard(PEChain_21_io_discard),
    .io_inData(PEChain_21_io_inData),
    .io_rightPropDiscard(PEChain_21_io_rightPropDiscard),
    .io_leftOutData(PEChain_21_io_leftOutData),
    .io_rightOutData(PEChain_21_io_rightOutData),
    .io_currDiscard(PEChain_21_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_21_io_toLeftPropDiscard)
  );
  PE_46 PEChain_22 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_22_clock),
    .reset(PEChain_22_reset),
    .io_enableSort(PEChain_22_io_enableSort),
    .io_state(PEChain_22_io_state),
    .io_leftNBR_data(PEChain_22_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_22_io_leftNBR_compRes),
    .io_rightNBR_data(PEChain_22_io_rightNBR_data),
    .io_rightNBR_compRes(PEChain_22_io_rightNBR_compRes),
    .io_currCell_data(PEChain_22_io_currCell_data),
    .io_currCell_compRes(PEChain_22_io_currCell_compRes),
    .io_lastCell(PEChain_22_io_lastCell),
    .io_active(PEChain_22_io_active),
    .io_discard(PEChain_22_io_discard),
    .io_inData(PEChain_22_io_inData),
    .io_rightPropDiscard(PEChain_22_io_rightPropDiscard),
    .io_leftOutData(PEChain_22_io_leftOutData),
    .io_rightOutData(PEChain_22_io_rightOutData),
    .io_currDiscard(PEChain_22_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_22_io_toLeftPropDiscard)
  );
  PE_47 PEChain_23 ( // @[LinearSorter.scala 143:24]
    .clock(PEChain_23_clock),
    .reset(PEChain_23_reset),
    .io_enableSort(PEChain_23_io_enableSort),
    .io_state(PEChain_23_io_state),
    .io_leftNBR_data(PEChain_23_io_leftNBR_data),
    .io_leftNBR_compRes(PEChain_23_io_leftNBR_compRes),
    .io_currCell_data(PEChain_23_io_currCell_data),
    .io_currCell_compRes(PEChain_23_io_currCell_compRes),
    .io_lastCell(PEChain_23_io_lastCell),
    .io_active(PEChain_23_io_active),
    .io_discard(PEChain_23_io_discard),
    .io_inData(PEChain_23_io_inData),
    .io_leftOutData(PEChain_23_io_leftOutData),
    .io_currDiscard(PEChain_23_io_currDiscard),
    .io_toLeftPropDiscard(PEChain_23_io_toLeftPropDiscard)
  );
  assign _T_1 = lisSizeReg - 6'h1; // @[LinearSorter.scala 86:43]
  assign _T_96 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_98 = cntInData + 5'h1; // @[LinearSorter.scala 92:28]
  assign _T_99 = state == 2'h0; // @[LinearSorter.scala 94:20]
  assign _GEN_111 = {{1'd0}, cntInData}; // @[LinearSorter.scala 98:19]
  assign _T_102 = _GEN_111 == _T_1; // @[LinearSorter.scala 98:19]
  assign _T_104 = _T_102 & _T_96; // @[LinearSorter.scala 98:42]
  assign _T_113 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_7 = _T_96 ? 2'h1 : state; // @[LinearSorter.scala 117:27]
  assign _T_115 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign fireLastIn = io_lastIn & _T_96; // @[LinearSorter.scala 111:30]
  assign _GEN_8 = fireLastIn ? 2'h2 : state; // @[LinearSorter.scala 120:62]
  assign _T_117 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_112 = {{1'd0}, cntOutData}; // @[LinearSorter.scala 125:28]
  assign _T_120 = _GEN_112 == _T_1; // @[LinearSorter.scala 125:28]
  assign _GEN_9 = _T_120 ? 2'h0 : state; // @[LinearSorter.scala 125:50]
  assign _GEN_10 = _T_117 ? _GEN_9 : state; // @[Conditional.scala 39:67]
  assign _GEN_11 = _T_115 ? _GEN_8 : _GEN_10; // @[Conditional.scala 39:67]
  assign state_next = _T_113 ? _GEN_7 : _GEN_11; // @[Conditional.scala 40:58]
  assign _T_105 = state_next == 2'h0; // @[LinearSorter.scala 101:25]
  assign _GEN_2 = _T_105 ? 1'h0 : initialInDone; // @[LinearSorter.scala 101:36]
  assign _GEN_3 = _T_104 | _GEN_2; // @[LinearSorter.scala 98:59]
  assign _T_106 = io_out_valid & io_out_ready; // @[LinearSorter.scala 106:29]
  assign _T_107 = state == 2'h2; // @[LinearSorter.scala 106:54]
  assign enable = _T_106 & _T_107; // @[LinearSorter.scala 106:45]
  assign _T_109 = cntOutData == 5'h17; // @[LISutil.scala 13:24]
  assign _T_111 = cntOutData + 5'h1; // @[LISutil.scala 14:22]
  assign _T_121 = state_next != 2'h2; // @[LinearSorter.scala 137:33]
  assign outputData_0 = PEChain_0_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign outputData_1 = PEChain_1_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_16 = 5'h1 == _T_1[4:0] ? $signed(outputData_1) : $signed(outputData_0); // @[LinearSorter.scala 137:21]
  assign outputData_2 = PEChain_2_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_17 = 5'h2 == _T_1[4:0] ? $signed(outputData_2) : $signed(_GEN_16); // @[LinearSorter.scala 137:21]
  assign outputData_3 = PEChain_3_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_18 = 5'h3 == _T_1[4:0] ? $signed(outputData_3) : $signed(_GEN_17); // @[LinearSorter.scala 137:21]
  assign outputData_4 = PEChain_4_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_19 = 5'h4 == _T_1[4:0] ? $signed(outputData_4) : $signed(_GEN_18); // @[LinearSorter.scala 137:21]
  assign outputData_5 = PEChain_5_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_20 = 5'h5 == _T_1[4:0] ? $signed(outputData_5) : $signed(_GEN_19); // @[LinearSorter.scala 137:21]
  assign outputData_6 = PEChain_6_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_21 = 5'h6 == _T_1[4:0] ? $signed(outputData_6) : $signed(_GEN_20); // @[LinearSorter.scala 137:21]
  assign outputData_7 = PEChain_7_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_22 = 5'h7 == _T_1[4:0] ? $signed(outputData_7) : $signed(_GEN_21); // @[LinearSorter.scala 137:21]
  assign outputData_8 = PEChain_8_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_23 = 5'h8 == _T_1[4:0] ? $signed(outputData_8) : $signed(_GEN_22); // @[LinearSorter.scala 137:21]
  assign outputData_9 = PEChain_9_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_24 = 5'h9 == _T_1[4:0] ? $signed(outputData_9) : $signed(_GEN_23); // @[LinearSorter.scala 137:21]
  assign outputData_10 = PEChain_10_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_25 = 5'ha == _T_1[4:0] ? $signed(outputData_10) : $signed(_GEN_24); // @[LinearSorter.scala 137:21]
  assign outputData_11 = PEChain_11_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_26 = 5'hb == _T_1[4:0] ? $signed(outputData_11) : $signed(_GEN_25); // @[LinearSorter.scala 137:21]
  assign outputData_12 = PEChain_12_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_27 = 5'hc == _T_1[4:0] ? $signed(outputData_12) : $signed(_GEN_26); // @[LinearSorter.scala 137:21]
  assign outputData_13 = PEChain_13_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_28 = 5'hd == _T_1[4:0] ? $signed(outputData_13) : $signed(_GEN_27); // @[LinearSorter.scala 137:21]
  assign outputData_14 = PEChain_14_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_29 = 5'he == _T_1[4:0] ? $signed(outputData_14) : $signed(_GEN_28); // @[LinearSorter.scala 137:21]
  assign outputData_15 = PEChain_15_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_30 = 5'hf == _T_1[4:0] ? $signed(outputData_15) : $signed(_GEN_29); // @[LinearSorter.scala 137:21]
  assign outputData_16 = PEChain_16_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_31 = 5'h10 == _T_1[4:0] ? $signed(outputData_16) : $signed(_GEN_30); // @[LinearSorter.scala 137:21]
  assign outputData_17 = PEChain_17_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_32 = 5'h11 == _T_1[4:0] ? $signed(outputData_17) : $signed(_GEN_31); // @[LinearSorter.scala 137:21]
  assign outputData_18 = PEChain_18_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_33 = 5'h12 == _T_1[4:0] ? $signed(outputData_18) : $signed(_GEN_32); // @[LinearSorter.scala 137:21]
  assign outputData_19 = PEChain_19_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_34 = 5'h13 == _T_1[4:0] ? $signed(outputData_19) : $signed(_GEN_33); // @[LinearSorter.scala 137:21]
  assign outputData_20 = PEChain_20_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_35 = 5'h14 == _T_1[4:0] ? $signed(outputData_20) : $signed(_GEN_34); // @[LinearSorter.scala 137:21]
  assign outputData_21 = PEChain_21_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_36 = 5'h15 == _T_1[4:0] ? $signed(outputData_21) : $signed(_GEN_35); // @[LinearSorter.scala 137:21]
  assign outputData_22 = PEChain_22_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_37 = 5'h16 == _T_1[4:0] ? $signed(outputData_22) : $signed(_GEN_36); // @[LinearSorter.scala 137:21]
  assign outputData_23 = PEChain_23_io_currCell_data; // @[LinearSorter.scala 73:24 LinearSorter.scala 170:23]
  assign _GEN_38 = 5'h17 == _T_1[4:0] ? $signed(outputData_23) : $signed(_GEN_37); // @[LinearSorter.scala 137:21]
  assign _T_136 = _T_107 & io_out_ready; // @[LinearSorter.scala 168:63]
  assign discardSignals_2 = PEChain_2_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_1 = PEChain_1_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_0 = PEChain_0_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_5 = PEChain_5_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_4 = PEChain_4_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_3 = PEChain_3_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_372 = {discardSignals_5,discardSignals_4,discardSignals_3,discardSignals_2,discardSignals_1,discardSignals_0}; // @[LinearSorter.scala 177:50]
  assign discardSignals_8 = PEChain_8_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_7 = PEChain_7_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_6 = PEChain_6_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_11 = PEChain_11_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_10 = PEChain_10_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_9 = PEChain_9_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_378 = {discardSignals_11,discardSignals_10,discardSignals_9,discardSignals_8,discardSignals_7,discardSignals_6,_T_372}; // @[LinearSorter.scala 177:50]
  assign discardSignals_14 = PEChain_14_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_13 = PEChain_13_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_12 = PEChain_12_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_17 = PEChain_17_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_16 = PEChain_16_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_15 = PEChain_15_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_383 = {discardSignals_17,discardSignals_16,discardSignals_15,discardSignals_14,discardSignals_13,discardSignals_12}; // @[LinearSorter.scala 177:50]
  assign discardSignals_20 = PEChain_20_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_19 = PEChain_19_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_18 = PEChain_18_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_23 = PEChain_23_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_22 = PEChain_22_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign discardSignals_21 = PEChain_21_io_currDiscard; // @[LinearSorter.scala 74:28 LinearSorter.scala 171:27]
  assign _T_390 = {discardSignals_23,discardSignals_22,discardSignals_21,discardSignals_20,discardSignals_19,discardSignals_18,_T_383,_T_378}; // @[LinearSorter.scala 177:50]
  assign _T_415 = _T_390[22] ? 5'h16 : 5'h17; // @[Mux.scala 47:69]
  assign _T_416 = _T_390[21] ? 5'h15 : _T_415; // @[Mux.scala 47:69]
  assign _T_417 = _T_390[20] ? 5'h14 : _T_416; // @[Mux.scala 47:69]
  assign _T_418 = _T_390[19] ? 5'h13 : _T_417; // @[Mux.scala 47:69]
  assign _T_419 = _T_390[18] ? 5'h12 : _T_418; // @[Mux.scala 47:69]
  assign _T_420 = _T_390[17] ? 5'h11 : _T_419; // @[Mux.scala 47:69]
  assign _T_421 = _T_390[16] ? 5'h10 : _T_420; // @[Mux.scala 47:69]
  assign _T_422 = _T_390[15] ? 5'hf : _T_421; // @[Mux.scala 47:69]
  assign _T_423 = _T_390[14] ? 5'he : _T_422; // @[Mux.scala 47:69]
  assign _T_424 = _T_390[13] ? 5'hd : _T_423; // @[Mux.scala 47:69]
  assign _T_425 = _T_390[12] ? 5'hc : _T_424; // @[Mux.scala 47:69]
  assign _T_426 = _T_390[11] ? 5'hb : _T_425; // @[Mux.scala 47:69]
  assign _T_427 = _T_390[10] ? 5'ha : _T_426; // @[Mux.scala 47:69]
  assign _T_428 = _T_390[9] ? 5'h9 : _T_427; // @[Mux.scala 47:69]
  assign _T_429 = _T_390[8] ? 5'h8 : _T_428; // @[Mux.scala 47:69]
  assign _T_430 = _T_390[7] ? 5'h7 : _T_429; // @[Mux.scala 47:69]
  assign _T_431 = _T_390[6] ? 5'h6 : _T_430; // @[Mux.scala 47:69]
  assign _T_432 = _T_390[5] ? 5'h5 : _T_431; // @[Mux.scala 47:69]
  assign _T_433 = _T_390[4] ? 5'h4 : _T_432; // @[Mux.scala 47:69]
  assign _T_434 = _T_390[3] ? 5'h3 : _T_433; // @[Mux.scala 47:69]
  assign _T_435 = _T_390[2] ? 5'h2 : _T_434; // @[Mux.scala 47:69]
  assign _T_436 = _T_390[1] ? 5'h1 : _T_435; // @[Mux.scala 47:69]
  assign getDiscarded = _T_390[0] ? 5'h0 : _T_436; // @[Mux.scala 47:69]
  assign _T_438 = state != 2'h2; // @[LinearSorter.scala 199:49]
  assign _GEN_88 = 5'h1 == getDiscarded ? $signed(outputData_1) : $signed(outputData_0); // @[LinearSorter.scala 206:15]
  assign _GEN_89 = 5'h2 == getDiscarded ? $signed(outputData_2) : $signed(_GEN_88); // @[LinearSorter.scala 206:15]
  assign _GEN_90 = 5'h3 == getDiscarded ? $signed(outputData_3) : $signed(_GEN_89); // @[LinearSorter.scala 206:15]
  assign _GEN_91 = 5'h4 == getDiscarded ? $signed(outputData_4) : $signed(_GEN_90); // @[LinearSorter.scala 206:15]
  assign _GEN_92 = 5'h5 == getDiscarded ? $signed(outputData_5) : $signed(_GEN_91); // @[LinearSorter.scala 206:15]
  assign _GEN_93 = 5'h6 == getDiscarded ? $signed(outputData_6) : $signed(_GEN_92); // @[LinearSorter.scala 206:15]
  assign _GEN_94 = 5'h7 == getDiscarded ? $signed(outputData_7) : $signed(_GEN_93); // @[LinearSorter.scala 206:15]
  assign _GEN_95 = 5'h8 == getDiscarded ? $signed(outputData_8) : $signed(_GEN_94); // @[LinearSorter.scala 206:15]
  assign _GEN_96 = 5'h9 == getDiscarded ? $signed(outputData_9) : $signed(_GEN_95); // @[LinearSorter.scala 206:15]
  assign _GEN_97 = 5'ha == getDiscarded ? $signed(outputData_10) : $signed(_GEN_96); // @[LinearSorter.scala 206:15]
  assign _GEN_98 = 5'hb == getDiscarded ? $signed(outputData_11) : $signed(_GEN_97); // @[LinearSorter.scala 206:15]
  assign _GEN_99 = 5'hc == getDiscarded ? $signed(outputData_12) : $signed(_GEN_98); // @[LinearSorter.scala 206:15]
  assign _GEN_100 = 5'hd == getDiscarded ? $signed(outputData_13) : $signed(_GEN_99); // @[LinearSorter.scala 206:15]
  assign _GEN_101 = 5'he == getDiscarded ? $signed(outputData_14) : $signed(_GEN_100); // @[LinearSorter.scala 206:15]
  assign _GEN_102 = 5'hf == getDiscarded ? $signed(outputData_15) : $signed(_GEN_101); // @[LinearSorter.scala 206:15]
  assign _GEN_103 = 5'h10 == getDiscarded ? $signed(outputData_16) : $signed(_GEN_102); // @[LinearSorter.scala 206:15]
  assign _GEN_104 = 5'h11 == getDiscarded ? $signed(outputData_17) : $signed(_GEN_103); // @[LinearSorter.scala 206:15]
  assign _GEN_105 = 5'h12 == getDiscarded ? $signed(outputData_18) : $signed(_GEN_104); // @[LinearSorter.scala 206:15]
  assign _GEN_106 = 5'h13 == getDiscarded ? $signed(outputData_19) : $signed(_GEN_105); // @[LinearSorter.scala 206:15]
  assign _GEN_107 = 5'h14 == getDiscarded ? $signed(outputData_20) : $signed(_GEN_106); // @[LinearSorter.scala 206:15]
  assign _GEN_108 = 5'h15 == getDiscarded ? $signed(outputData_21) : $signed(_GEN_107); // @[LinearSorter.scala 206:15]
  assign _GEN_109 = 5'h16 == getDiscarded ? $signed(outputData_22) : $signed(_GEN_108); // @[LinearSorter.scala 206:15]
  assign _T_444 = ~initialInDone; // @[LinearSorter.scala 208:18]
  assign _T_446 = io_out_ready & _T_438; // @[LinearSorter.scala 208:49]
  assign _T_448 = initialInDone & io_in_valid; // @[LinearSorter.scala 209:33]
  assign io_in_ready = _T_444 | _T_446; // @[LinearSorter.scala 208:15]
  assign io_out_valid = _T_448 | _T_107; // @[LinearSorter.scala 209:16]
  assign io_out_bits = 5'h17 == getDiscarded ? $signed(outputData_23) : $signed(_GEN_109); // @[LinearSorter.scala 206:15]
  assign io_lastOut = _GEN_112 == _T_1; // @[LinearSorter.scala 207:15]
  assign io_sortedData_0 = PEChain_0_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_1 = PEChain_1_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_2 = PEChain_2_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_3 = PEChain_3_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_4 = PEChain_4_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_5 = PEChain_5_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_6 = PEChain_6_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_7 = PEChain_7_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_8 = PEChain_8_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_9 = PEChain_9_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_10 = PEChain_10_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_11 = PEChain_11_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_12 = PEChain_12_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_13 = PEChain_13_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_14 = PEChain_14_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_15 = PEChain_15_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_16 = PEChain_16_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_17 = PEChain_17_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_18 = PEChain_18_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_19 = PEChain_19_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_20 = PEChain_20_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_21 = PEChain_21_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_22 = PEChain_22_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sortedData_23 = PEChain_23_io_currCell_data; // @[LinearSorter.scala 205:17]
  assign io_sorterFull = initialInDone & _T_438; // @[LinearSorter.scala 199:23]
  assign io_sorterEmpty = state == 2'h0; // @[LinearSorter.scala 202:24]
  assign PEChain_0_clock = clock;
  assign PEChain_0_reset = reset;
  assign PEChain_0_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_0_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_0_io_rightNBR_data = PEChain_1_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_0_io_rightNBR_compRes = PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_0_io_lastCell = 6'h0 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_0_io_discard = _T_107 & initialInDone; // @[LinearSorter.scala 156:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_0_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_0_io_rightPropDiscard = PEChain_1_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_1_clock = clock;
  assign PEChain_1_reset = reset;
  assign PEChain_1_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_1_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_1_io_leftNBR_data = PEChain_0_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_1_io_leftNBR_compRes = PEChain_0_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_1_io_rightNBR_data = PEChain_2_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_1_io_rightNBR_compRes = PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_1_io_lastCell = 6'h1 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_1_io_active = 6'h1 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_1_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_1_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_1_io_rightPropDiscard = PEChain_2_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_2_clock = clock;
  assign PEChain_2_reset = reset;
  assign PEChain_2_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_2_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_2_io_leftNBR_data = PEChain_1_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_2_io_leftNBR_compRes = PEChain_1_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_2_io_rightNBR_data = PEChain_3_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_2_io_rightNBR_compRes = PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_2_io_lastCell = 6'h2 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_2_io_active = 6'h2 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_2_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_2_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_2_io_rightPropDiscard = PEChain_3_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_3_clock = clock;
  assign PEChain_3_reset = reset;
  assign PEChain_3_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_3_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_3_io_leftNBR_data = PEChain_2_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_3_io_leftNBR_compRes = PEChain_2_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_3_io_rightNBR_data = PEChain_4_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_3_io_rightNBR_compRes = PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_3_io_lastCell = 6'h3 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_3_io_active = 6'h3 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_3_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_3_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_3_io_rightPropDiscard = PEChain_4_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_4_clock = clock;
  assign PEChain_4_reset = reset;
  assign PEChain_4_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_4_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_4_io_leftNBR_data = PEChain_3_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_4_io_leftNBR_compRes = PEChain_3_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_4_io_rightNBR_data = PEChain_5_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_4_io_rightNBR_compRes = PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_4_io_lastCell = 6'h4 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_4_io_active = 6'h4 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_4_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_4_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_4_io_rightPropDiscard = PEChain_5_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_5_clock = clock;
  assign PEChain_5_reset = reset;
  assign PEChain_5_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_5_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_5_io_leftNBR_data = PEChain_4_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_5_io_leftNBR_compRes = PEChain_4_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_5_io_rightNBR_data = PEChain_6_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_5_io_rightNBR_compRes = PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_5_io_lastCell = 6'h5 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_5_io_active = 6'h5 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_5_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_5_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_5_io_rightPropDiscard = PEChain_6_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_6_clock = clock;
  assign PEChain_6_reset = reset;
  assign PEChain_6_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_6_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_6_io_leftNBR_data = PEChain_5_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_6_io_leftNBR_compRes = PEChain_5_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_6_io_rightNBR_data = PEChain_7_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_6_io_rightNBR_compRes = PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_6_io_lastCell = 6'h6 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_6_io_active = 6'h6 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_6_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_6_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_6_io_rightPropDiscard = PEChain_7_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_7_clock = clock;
  assign PEChain_7_reset = reset;
  assign PEChain_7_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_7_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_7_io_leftNBR_data = PEChain_6_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_7_io_leftNBR_compRes = PEChain_6_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_7_io_rightNBR_data = PEChain_8_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_7_io_rightNBR_compRes = PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_7_io_lastCell = 6'h7 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_7_io_active = 6'h7 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_7_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_7_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_7_io_rightPropDiscard = PEChain_8_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_8_clock = clock;
  assign PEChain_8_reset = reset;
  assign PEChain_8_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_8_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_8_io_leftNBR_data = PEChain_7_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_8_io_leftNBR_compRes = PEChain_7_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_8_io_rightNBR_data = PEChain_9_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_8_io_rightNBR_compRes = PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_8_io_lastCell = 6'h8 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_8_io_active = 6'h8 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_8_io_discard = _T_107 ? 1'h0 : initialInDone; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_8_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_8_io_rightPropDiscard = PEChain_9_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_9_clock = clock;
  assign PEChain_9_reset = reset;
  assign PEChain_9_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_9_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_9_io_leftNBR_data = PEChain_8_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_9_io_leftNBR_compRes = PEChain_8_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_9_io_rightNBR_data = PEChain_10_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_9_io_rightNBR_compRes = PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_9_io_lastCell = 6'h9 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_9_io_active = 6'h9 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_9_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_9_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_9_io_rightPropDiscard = PEChain_10_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_10_clock = clock;
  assign PEChain_10_reset = reset;
  assign PEChain_10_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_10_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_10_io_leftNBR_data = PEChain_9_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_10_io_leftNBR_compRes = PEChain_9_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_10_io_rightNBR_data = PEChain_11_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_10_io_rightNBR_compRes = PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_10_io_lastCell = 6'ha == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_10_io_active = 6'ha <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_10_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_10_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_10_io_rightPropDiscard = PEChain_11_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_11_clock = clock;
  assign PEChain_11_reset = reset;
  assign PEChain_11_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_11_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_11_io_leftNBR_data = PEChain_10_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_11_io_leftNBR_compRes = PEChain_10_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_11_io_rightNBR_data = PEChain_12_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_11_io_rightNBR_compRes = PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_11_io_lastCell = 6'hb == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_11_io_active = 6'hb <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_11_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_11_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_11_io_rightPropDiscard = PEChain_12_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_12_clock = clock;
  assign PEChain_12_reset = reset;
  assign PEChain_12_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_12_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_12_io_leftNBR_data = PEChain_11_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_12_io_leftNBR_compRes = PEChain_11_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_12_io_rightNBR_data = PEChain_13_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_12_io_rightNBR_compRes = PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_12_io_lastCell = 6'hc == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_12_io_active = 6'hc <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_12_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_12_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_12_io_rightPropDiscard = PEChain_13_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_13_clock = clock;
  assign PEChain_13_reset = reset;
  assign PEChain_13_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_13_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_13_io_leftNBR_data = PEChain_12_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_13_io_leftNBR_compRes = PEChain_12_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_13_io_rightNBR_data = PEChain_14_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_13_io_rightNBR_compRes = PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_13_io_lastCell = 6'hd == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_13_io_active = 6'hd <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_13_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_13_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_13_io_rightPropDiscard = PEChain_14_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_14_clock = clock;
  assign PEChain_14_reset = reset;
  assign PEChain_14_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_14_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_14_io_leftNBR_data = PEChain_13_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_14_io_leftNBR_compRes = PEChain_13_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_14_io_rightNBR_data = PEChain_15_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_14_io_rightNBR_compRes = PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_14_io_lastCell = 6'he == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_14_io_active = 6'he <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_14_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_14_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_14_io_rightPropDiscard = PEChain_15_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_15_clock = clock;
  assign PEChain_15_reset = reset;
  assign PEChain_15_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_15_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_15_io_leftNBR_data = PEChain_14_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_15_io_leftNBR_compRes = PEChain_14_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_15_io_rightNBR_data = PEChain_16_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_15_io_rightNBR_compRes = PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_15_io_lastCell = 6'hf == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_15_io_active = 6'hf <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_15_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_15_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_15_io_rightPropDiscard = PEChain_16_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_16_clock = clock;
  assign PEChain_16_reset = reset;
  assign PEChain_16_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_16_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_16_io_leftNBR_data = PEChain_15_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_16_io_leftNBR_compRes = PEChain_15_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_16_io_rightNBR_data = PEChain_17_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_16_io_rightNBR_compRes = PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_16_io_lastCell = 6'h10 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_16_io_active = 6'h10 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_16_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_16_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_16_io_rightPropDiscard = PEChain_17_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_17_clock = clock;
  assign PEChain_17_reset = reset;
  assign PEChain_17_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_17_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_17_io_leftNBR_data = PEChain_16_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_17_io_leftNBR_compRes = PEChain_16_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_17_io_rightNBR_data = PEChain_18_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_17_io_rightNBR_compRes = PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_17_io_lastCell = 6'h11 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_17_io_active = 6'h11 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_17_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_17_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_17_io_rightPropDiscard = PEChain_18_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_18_clock = clock;
  assign PEChain_18_reset = reset;
  assign PEChain_18_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_18_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_18_io_leftNBR_data = PEChain_17_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_18_io_leftNBR_compRes = PEChain_17_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_18_io_rightNBR_data = PEChain_19_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_18_io_rightNBR_compRes = PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_18_io_lastCell = 6'h12 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_18_io_active = 6'h12 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_18_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_18_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_18_io_rightPropDiscard = PEChain_19_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_19_clock = clock;
  assign PEChain_19_reset = reset;
  assign PEChain_19_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_19_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_19_io_leftNBR_data = PEChain_18_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_19_io_leftNBR_compRes = PEChain_18_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_19_io_rightNBR_data = PEChain_20_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_19_io_rightNBR_compRes = PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_19_io_lastCell = 6'h13 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_19_io_active = 6'h13 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_19_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_19_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_19_io_rightPropDiscard = PEChain_20_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_20_clock = clock;
  assign PEChain_20_reset = reset;
  assign PEChain_20_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_20_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_20_io_leftNBR_data = PEChain_19_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_20_io_leftNBR_compRes = PEChain_19_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_20_io_rightNBR_data = PEChain_21_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_20_io_rightNBR_compRes = PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_20_io_lastCell = 6'h14 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_20_io_active = 6'h14 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_20_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_20_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_20_io_rightPropDiscard = PEChain_21_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_21_clock = clock;
  assign PEChain_21_reset = reset;
  assign PEChain_21_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_21_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_21_io_leftNBR_data = PEChain_20_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_21_io_leftNBR_compRes = PEChain_20_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_21_io_rightNBR_data = PEChain_22_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_21_io_rightNBR_compRes = PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_21_io_lastCell = 6'h15 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_21_io_active = 6'h15 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_21_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_21_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_21_io_rightPropDiscard = PEChain_22_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_22_clock = clock;
  assign PEChain_22_reset = reset;
  assign PEChain_22_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_22_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_22_io_leftNBR_data = PEChain_21_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_22_io_leftNBR_compRes = PEChain_21_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_22_io_rightNBR_data = PEChain_23_io_leftOutData; // @[LinearSorter.scala 190:30]
  assign PEChain_22_io_rightNBR_compRes = PEChain_23_io_currCell_compRes; // @[LinearSorter.scala 191:33]
  assign PEChain_22_io_lastCell = 6'h16 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_22_io_active = 6'h16 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_22_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_22_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
  assign PEChain_22_io_rightPropDiscard = PEChain_23_io_toLeftPropDiscard; // @[LinearSorter.scala 193:34]
  assign PEChain_23_clock = clock;
  assign PEChain_23_reset = reset;
  assign PEChain_23_io_enableSort = _T_96 | _T_136; // @[LinearSorter.scala 168:26]
  assign PEChain_23_io_state = _T_113 ? _GEN_7 : _GEN_11; // @[LinearSorter.scala 169:21]
  assign PEChain_23_io_leftNBR_data = PEChain_22_io_rightOutData; // @[LinearSorter.scala 187:29]
  assign PEChain_23_io_leftNBR_compRes = PEChain_22_io_currCell_compRes; // @[LinearSorter.scala 188:32]
  assign PEChain_23_io_lastCell = 6'h17 == _T_1; // @[LinearSorter.scala 148:30]
  assign PEChain_23_io_active = 6'h17 <= _T_1; // @[LinearSorter.scala 147:28]
  assign PEChain_23_io_discard = 1'h0; // @[LinearSorter.scala 158:33 LinearSorter.scala 161:31 LinearSorter.scala 164:31]
  assign PEChain_23_io_inData = _T_121 ? $signed(io_in_bits) : $signed(_GEN_38); // @[LinearSorter.scala 144:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  initialInDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cntInData = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  lisSizeReg = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cntOutData = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      initialInDone <= 1'h0;
    end else begin
      initialInDone <= _GEN_3;
    end
    if (reset) begin
      cntInData <= 5'h0;
    end else if (_T_96) begin
      cntInData <= _T_98;
    end else if (_T_99) begin
      cntInData <= 5'h0;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_113) begin
      if (_T_96) begin
        state <= 2'h1;
      end
    end else if (_T_115) begin
      if (fireLastIn) begin
        state <= 2'h2;
      end
    end else if (_T_117) begin
      if (_T_120) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      lisSizeReg <= 6'h18;
    end else if (_T_113) begin
      lisSizeReg <= io_lisSize;
    end
    if (reset) begin
      cntOutData <= 5'h0;
    end else if (_T_99) begin
      cntOutData <= 5'h0;
    end else if (enable) begin
      if (_T_109) begin
        cntOutData <= 5'h0;
      end else begin
        cntOutData <= _T_111;
      end
    end
  end
endmodule
module AXI4LISBlock_2(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  lis_clock; // @[LISDspBlock.scala 55:21]
  wire  lis_reset; // @[LISDspBlock.scala 55:21]
  wire  lis_io_in_ready; // @[LISDspBlock.scala 55:21]
  wire  lis_io_in_valid; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_in_bits; // @[LISDspBlock.scala 55:21]
  wire  lis_io_lastIn; // @[LISDspBlock.scala 55:21]
  wire  lis_io_out_ready; // @[LISDspBlock.scala 55:21]
  wire  lis_io_out_valid; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_out_bits; // @[LISDspBlock.scala 55:21]
  wire  lis_io_lastOut; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_0; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_1; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_2; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_3; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_4; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_5; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_6; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_7; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_8; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_9; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_10; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_11; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_12; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_13; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_14; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_15; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_16; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_17; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_18; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_19; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_20; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_21; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_22; // @[LISDspBlock.scala 55:21]
  wire [15:0] lis_io_sortedData_23; // @[LISDspBlock.scala 55:21]
  wire  lis_io_sorterFull; // @[LISDspBlock.scala 55:21]
  wire  lis_io_sorterEmpty; // @[LISDspBlock.scala 55:21]
  wire [5:0] lis_io_lisSize; // @[LISDspBlock.scala 55:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  sortDir; // @[LISDspBlock.scala 58:26]
  reg [31:0] _RAND_0;
  reg  flushData; // @[LISDspBlock.scala 59:28]
  reg [31:0] _RAND_1;
  reg [4:0] discardPos; // @[LISDspBlock.scala 60:29]
  reg [31:0] _RAND_2;
  reg [4:0] sendOnOutput; // @[LISDspBlock.scala 61:31]
  reg [31:0] _RAND_3;
  reg [4:0] lisSize; // @[LISDspBlock.scala 62:26]
  reg [31:0] _RAND_4;
  reg  sorterFull; // @[LISDspBlock.scala 65:29]
  reg [31:0] _RAND_5;
  reg  sorterEmpty; // @[LISDspBlock.scala 66:30]
  reg [31:0] _RAND_6;
  wire [31:0] _T_2; // @[LISDspBlock.scala 71:44]
  wire [15:0] _GEN_0; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_1; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_2; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_3; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_4; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_5; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_6; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_7; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_8; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_9; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_10; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_11; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_12; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_13; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_14; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_15; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_16; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_17; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_18; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_19; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_20; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_21; // @[LISDspBlock.scala 92:82]
  wire [15:0] _GEN_22; // @[LISDspBlock.scala 92:82]
  wire [15:0] _T_4; // @[LISDspBlock.scala 92:82]
  wire  _T_7; // @[RegisterRouter.scala 40:39]
  wire  _T_8; // @[RegisterRouter.scala 40:26]
  wire  _T_9; // @[RegisterRouter.scala 42:29]
  wire  _T_52_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_16; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_281; // @[Cat.scala 29:58]
  wire [5:0] _T_56; // @[RegisterRouter.scala 59:16]
  wire  _T_64; // @[RegisterRouter.scala 59:16]
  wire  _T_10; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_19; // @[OneHot.scala 65:12]
  wire [1:0] _T_21; // @[Misc.scala 200:81]
  wire  _T_22; // @[Misc.scala 204:21]
  wire  _T_25; // @[Misc.scala 209:20]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_30; // @[Misc.scala 213:38]
  wire  _T_31; // @[Misc.scala 213:29]
  wire  _T_34; // @[Misc.scala 209:20]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire  _T_44; // @[Misc.scala 212:27]
  wire  _T_45; // @[Misc.scala 213:38]
  wire  _T_46; // @[Misc.scala 213:29]
  wire [3:0] _T_49; // @[Cat.scala 29:58]
  wire [3:0] _T_51; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_80; // @[Bitwise.scala 72:12]
  wire [7:0] _T_82; // @[Bitwise.scala 72:12]
  wire [7:0] _T_84; // @[Bitwise.scala 72:12]
  wire [7:0] _T_86; // @[Bitwise.scala 72:12]
  wire [31:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_300; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_282; // @[OneHot.scala 58:35]
  wire  _T_347; // @[RegisterRouter.scala 59:16]
  wire  _T_349; // @[RegisterRouter.scala 59:16]
  wire  _T_350; // @[RegisterRouter.scala 59:16]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _GEN_24; // @[RegField.scala 134:88]
  wire  _T_154; // @[RegisterRouter.scala 59:16]
  wire  _T_354; // @[RegisterRouter.scala 59:16]
  wire  _T_355; // @[RegisterRouter.scala 59:16]
  wire  _T_161; // @[RegisterRouter.scala 59:16]
  wire  _T_359; // @[RegisterRouter.scala 59:16]
  wire  _T_360; // @[RegisterRouter.scala 59:16]
  wire  _T_207; // @[RegisterRouter.scala 59:16]
  wire  _T_364; // @[RegisterRouter.scala 59:16]
  wire  _T_365; // @[RegisterRouter.scala 59:16]
  wire  _T_230; // @[RegisterRouter.scala 59:16]
  wire  _T_369; // @[RegisterRouter.scala 59:16]
  wire  _T_370; // @[RegisterRouter.scala 59:16]
  wire  _T_253; // @[RegisterRouter.scala 59:16]
  wire  _GEN_62; // @[MuxLiteral.scala 48:10]
  wire  _GEN_63; // @[MuxLiteral.scala 48:10]
  wire  _GEN_64; // @[MuxLiteral.scala 48:10]
  wire  _GEN_65; // @[MuxLiteral.scala 48:10]
  wire  _GEN_66; // @[MuxLiteral.scala 48:10]
  wire  _GEN_67; // @[MuxLiteral.scala 48:10]
  wire  _GEN_77; // @[MuxLiteral.scala 48:10]
  wire  _GEN_68; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_0; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_70; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_71; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_72; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_73; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_74; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_492_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [4:0] _GEN_75; // @[MuxLiteral.scala 48:10]
  wire [4:0] _GEN_76; // @[MuxLiteral.scala 48:10]
  wire [4:0] _T_494; // @[RegisterRouter.scala 59:16]
  wire  _T_495_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_495_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_498; // @[RegisterRouter.scala 65:29]
  LinearSorter_2 lis ( // @[LISDspBlock.scala 55:21]
    .clock(lis_clock),
    .reset(lis_reset),
    .io_in_ready(lis_io_in_ready),
    .io_in_valid(lis_io_in_valid),
    .io_in_bits(lis_io_in_bits),
    .io_lastIn(lis_io_lastIn),
    .io_out_ready(lis_io_out_ready),
    .io_out_valid(lis_io_out_valid),
    .io_out_bits(lis_io_out_bits),
    .io_lastOut(lis_io_lastOut),
    .io_sortedData_0(lis_io_sortedData_0),
    .io_sortedData_1(lis_io_sortedData_1),
    .io_sortedData_2(lis_io_sortedData_2),
    .io_sortedData_3(lis_io_sortedData_3),
    .io_sortedData_4(lis_io_sortedData_4),
    .io_sortedData_5(lis_io_sortedData_5),
    .io_sortedData_6(lis_io_sortedData_6),
    .io_sortedData_7(lis_io_sortedData_7),
    .io_sortedData_8(lis_io_sortedData_8),
    .io_sortedData_9(lis_io_sortedData_9),
    .io_sortedData_10(lis_io_sortedData_10),
    .io_sortedData_11(lis_io_sortedData_11),
    .io_sortedData_12(lis_io_sortedData_12),
    .io_sortedData_13(lis_io_sortedData_13),
    .io_sortedData_14(lis_io_sortedData_14),
    .io_sortedData_15(lis_io_sortedData_15),
    .io_sortedData_16(lis_io_sortedData_16),
    .io_sortedData_17(lis_io_sortedData_17),
    .io_sortedData_18(lis_io_sortedData_18),
    .io_sortedData_19(lis_io_sortedData_19),
    .io_sortedData_20(lis_io_sortedData_20),
    .io_sortedData_21(lis_io_sortedData_21),
    .io_sortedData_22(lis_io_sortedData_22),
    .io_sortedData_23(lis_io_sortedData_23),
    .io_sorterFull(lis_io_sorterFull),
    .io_sorterEmpty(lis_io_sorterEmpty),
    .io_lisSize(lis_io_lisSize)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_2 = auto_stream_in_bits_data; // @[LISDspBlock.scala 71:44]
  assign _GEN_0 = lis_io_sortedData_0; // @[LISDspBlock.scala 92:82]
  assign _GEN_1 = 5'h1 == sendOnOutput ? $signed(lis_io_sortedData_1) : $signed(_GEN_0); // @[LISDspBlock.scala 92:82]
  assign _GEN_2 = 5'h2 == sendOnOutput ? $signed(lis_io_sortedData_2) : $signed(_GEN_1); // @[LISDspBlock.scala 92:82]
  assign _GEN_3 = 5'h3 == sendOnOutput ? $signed(lis_io_sortedData_3) : $signed(_GEN_2); // @[LISDspBlock.scala 92:82]
  assign _GEN_4 = 5'h4 == sendOnOutput ? $signed(lis_io_sortedData_4) : $signed(_GEN_3); // @[LISDspBlock.scala 92:82]
  assign _GEN_5 = 5'h5 == sendOnOutput ? $signed(lis_io_sortedData_5) : $signed(_GEN_4); // @[LISDspBlock.scala 92:82]
  assign _GEN_6 = 5'h6 == sendOnOutput ? $signed(lis_io_sortedData_6) : $signed(_GEN_5); // @[LISDspBlock.scala 92:82]
  assign _GEN_7 = 5'h7 == sendOnOutput ? $signed(lis_io_sortedData_7) : $signed(_GEN_6); // @[LISDspBlock.scala 92:82]
  assign _GEN_8 = 5'h8 == sendOnOutput ? $signed(lis_io_sortedData_8) : $signed(_GEN_7); // @[LISDspBlock.scala 92:82]
  assign _GEN_9 = 5'h9 == sendOnOutput ? $signed(lis_io_sortedData_9) : $signed(_GEN_8); // @[LISDspBlock.scala 92:82]
  assign _GEN_10 = 5'ha == sendOnOutput ? $signed(lis_io_sortedData_10) : $signed(_GEN_9); // @[LISDspBlock.scala 92:82]
  assign _GEN_11 = 5'hb == sendOnOutput ? $signed(lis_io_sortedData_11) : $signed(_GEN_10); // @[LISDspBlock.scala 92:82]
  assign _GEN_12 = 5'hc == sendOnOutput ? $signed(lis_io_sortedData_12) : $signed(_GEN_11); // @[LISDspBlock.scala 92:82]
  assign _GEN_13 = 5'hd == sendOnOutput ? $signed(lis_io_sortedData_13) : $signed(_GEN_12); // @[LISDspBlock.scala 92:82]
  assign _GEN_14 = 5'he == sendOnOutput ? $signed(lis_io_sortedData_14) : $signed(_GEN_13); // @[LISDspBlock.scala 92:82]
  assign _GEN_15 = 5'hf == sendOnOutput ? $signed(lis_io_sortedData_15) : $signed(_GEN_14); // @[LISDspBlock.scala 92:82]
  assign _GEN_16 = 5'h10 == sendOnOutput ? $signed(lis_io_sortedData_16) : $signed(_GEN_15); // @[LISDspBlock.scala 92:82]
  assign _GEN_17 = 5'h11 == sendOnOutput ? $signed(lis_io_sortedData_17) : $signed(_GEN_16); // @[LISDspBlock.scala 92:82]
  assign _GEN_18 = 5'h12 == sendOnOutput ? $signed(lis_io_sortedData_18) : $signed(_GEN_17); // @[LISDspBlock.scala 92:82]
  assign _GEN_19 = 5'h13 == sendOnOutput ? $signed(lis_io_sortedData_19) : $signed(_GEN_18); // @[LISDspBlock.scala 92:82]
  assign _GEN_20 = 5'h14 == sendOnOutput ? $signed(lis_io_sortedData_20) : $signed(_GEN_19); // @[LISDspBlock.scala 92:82]
  assign _GEN_21 = 5'h15 == sendOnOutput ? $signed(lis_io_sortedData_21) : $signed(_GEN_20); // @[LISDspBlock.scala 92:82]
  assign _GEN_22 = 5'h16 == sendOnOutput ? $signed(lis_io_sortedData_22) : $signed(_GEN_21); // @[LISDspBlock.scala 92:82]
  assign _T_4 = 5'h17 == sendOnOutput ? $signed(lis_io_sortedData_23) : $signed(_GEN_22); // @[LISDspBlock.scala 92:82]
  assign _T_7 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_8 = auto_mem_in_ar_valid | _T_7; // @[RegisterRouter.scala 40:26]
  assign _T_9 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_52_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_16 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_281 = {_T_16[4],_T_16[3],_T_16[2]}; // @[Cat.scala 29:58]
  assign _T_56 = _T_16[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_64 = _T_56 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_10 = _T_52_ready & _T_9; // @[RegisterRouter.scala 42:26]
  assign _T_19 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_21 = _T_19 | 2'h1; // @[Misc.scala 200:81]
  assign _T_22 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_25 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_27 = _T_21[1] & _T_25; // @[Misc.scala 213:38]
  assign _T_28 = _T_22 | _T_27; // @[Misc.scala 213:29]
  assign _T_30 = _T_21[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_31 = _T_22 | _T_30; // @[Misc.scala 213:29]
  assign _T_34 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_35 = _T_25 & _T_34; // @[Misc.scala 212:27]
  assign _T_36 = _T_21[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_28 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = _T_25 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_39 = _T_21[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & _T_34; // @[Misc.scala 212:27]
  assign _T_42 = _T_21[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_31 | _T_42; // @[Misc.scala 213:29]
  assign _T_44 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_45 = _T_21[0] & _T_44; // @[Misc.scala 213:38]
  assign _T_46 = _T_31 | _T_45; // @[Misc.scala 213:29]
  assign _T_49 = {_T_46,_T_43,_T_40,_T_37}; // @[Cat.scala 29:58]
  assign _T_51 = auto_mem_in_ar_valid ? _T_49 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_80 = _T_51[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_82 = _T_51[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_84 = _T_51[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_86 = _T_51[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = {_T_86,_T_84,_T_82,_T_80}; // @[Cat.scala 29:58]
  assign _T_300 = _T_8 & _T_52_ready; // @[RegisterRouter.scala 59:16]
  assign _T_282 = 8'h1 << _T_281; // @[OneHot.scala 58:35]
  assign _T_347 = _T_300 & _T_9; // @[RegisterRouter.scala 59:16]
  assign _T_349 = _T_347 & _T_282[0]; // @[RegisterRouter.scala 59:16]
  assign _T_350 = _T_349 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_115 = _T_350 & _T_89[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_24 = _T_115 ? auto_mem_in_w_bits_data[0] : sortDir; // @[RegField.scala 134:88]
  assign _T_154 = _T_89[4:0] == 5'h1f; // @[RegisterRouter.scala 59:16]
  assign _T_354 = _T_347 & _T_282[1]; // @[RegisterRouter.scala 59:16]
  assign _T_355 = _T_354 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_161 = _T_355 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _T_359 = _T_347 & _T_282[2]; // @[RegisterRouter.scala 59:16]
  assign _T_360 = _T_359 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_207 = _T_360 & _T_89[0]; // @[RegisterRouter.scala 59:16]
  assign _T_364 = _T_347 & _T_282[3]; // @[RegisterRouter.scala 59:16]
  assign _T_365 = _T_364 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_230 = _T_365 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _T_369 = _T_347 & _T_282[4]; // @[RegisterRouter.scala 59:16]
  assign _T_370 = _T_369 & _T_64; // @[RegisterRouter.scala 59:16]
  assign _T_253 = _T_370 & _T_154; // @[RegisterRouter.scala 59:16]
  assign _GEN_62 = 3'h1 == _T_281 ? _T_64 : _T_64; // @[MuxLiteral.scala 48:10]
  assign _GEN_63 = 3'h2 == _T_281 ? _T_64 : _GEN_62; // @[MuxLiteral.scala 48:10]
  assign _GEN_64 = 3'h3 == _T_281 ? _T_64 : _GEN_63; // @[MuxLiteral.scala 48:10]
  assign _GEN_65 = 3'h4 == _T_281 ? _T_64 : _GEN_64; // @[MuxLiteral.scala 48:10]
  assign _GEN_66 = 3'h5 == _T_281 ? _T_64 : _GEN_65; // @[MuxLiteral.scala 48:10]
  assign _GEN_67 = 3'h6 == _T_281 ? _T_64 : _GEN_66; // @[MuxLiteral.scala 48:10]
  assign _GEN_77 = 3'h7 == _T_281; // @[MuxLiteral.scala 48:10]
  assign _GEN_68 = _GEN_77 | _GEN_67; // @[MuxLiteral.scala 48:10]
  assign _T_492_0 = {{4'd0}, sortDir}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_70 = 3'h1 == _T_281 ? lisSize : _T_492_0; // @[MuxLiteral.scala 48:10]
  assign _T_492_2 = {{4'd0}, flushData}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_71 = 3'h2 == _T_281 ? _T_492_2 : _GEN_70; // @[MuxLiteral.scala 48:10]
  assign _GEN_72 = 3'h3 == _T_281 ? discardPos : _GEN_71; // @[MuxLiteral.scala 48:10]
  assign _GEN_73 = 3'h4 == _T_281 ? sendOnOutput : _GEN_72; // @[MuxLiteral.scala 48:10]
  assign _T_492_5 = {{4'd0}, sorterFull}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_74 = 3'h5 == _T_281 ? _T_492_5 : _GEN_73; // @[MuxLiteral.scala 48:10]
  assign _T_492_6 = {{4'd0}, sorterEmpty}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_75 = 3'h6 == _T_281 ? _T_492_6 : _GEN_74; // @[MuxLiteral.scala 48:10]
  assign _GEN_76 = 3'h7 == _T_281 ? 5'h0 : _GEN_75; // @[MuxLiteral.scala 48:10]
  assign _T_494 = _GEN_68 ? _GEN_76 : 5'h0; // @[RegisterRouter.scala 59:16]
  assign _T_495_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_495_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_498 = ~_T_495_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_10 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_10 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_495_valid & _T_498; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_495_valid & _T_495_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = lis_io_in_ready; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = lis_io_out_valid; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {lis_io_out_bits,_T_4}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = lis_io_lastOut; // @[LazyModule.scala 173:49]
  assign lis_clock = clock;
  assign lis_reset = reset;
  assign lis_io_in_valid = auto_stream_in_valid; // @[LISDspBlock.scala 70:21]
  assign lis_io_in_bits = _T_2[15:0]; // @[LISDspBlock.scala 71:20]
  assign lis_io_lastIn = auto_stream_in_bits_last; // @[LISDspBlock.scala 69:19]
  assign lis_io_out_ready = auto_stream_out_ready; // @[LISDspBlock.scala 91:22]
  assign lis_io_lisSize = {{1'd0}, lisSize}; // @[LISDspBlock.scala 79:26]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_7; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{27'd0}, _T_494}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_495_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sortDir = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  flushData = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  discardPos = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sendOnOutput = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  lisSize = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sorterFull = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sorterEmpty = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    sortDir <= reset | _GEN_24;
    if (reset) begin
      flushData <= 1'h0;
    end else if (_T_207) begin
      flushData <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      discardPos <= 5'h0;
    end else if (_T_230) begin
      discardPos <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      sendOnOutput <= 5'h0;
    end else if (_T_253) begin
      sendOnOutput <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      lisSize <= 5'h18;
    end else if (_T_161) begin
      lisSize <= auto_mem_in_w_bits_data[4:0];
    end
    if (reset) begin
      sorterFull <= 1'h0;
    end else begin
      sorterFull <= lis_io_sorterFull;
    end
    sorterEmpty <= reset | lis_io_sorterEmpty;
  end
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  input   io_increment,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4,
  output  io_out_5,
  output  io_out_6,
  output  io_out_7,
  output  io_out_8,
  output  io_out_9,
  output  io_out_10,
  output  io_out_11,
  output  io_out_12,
  output  io_out_13,
  output  io_out_14,
  output  io_out_15
);
  reg  state_0; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_0;
  reg  state_1; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_1;
  reg  state_2; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_2;
  reg  state_3; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_3;
  reg  state_4; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_4;
  reg  state_5; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_5;
  reg  state_6; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_6;
  reg  state_7; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_7;
  reg  state_8; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_8;
  reg  state_9; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_9;
  reg  state_10; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_10;
  reg  state_11; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_11;
  reg  state_12; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_12;
  reg  state_13; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_13;
  reg  state_14; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_14;
  reg  state_15; // @[PRNG.scala 47:50]
  reg [31:0] _RAND_15;
  wire  _T_1; // @[LFSR.scala 15:41]
  wire  _T_2; // @[LFSR.scala 15:41]
  wire  _T_3; // @[LFSR.scala 15:41]
  wire  _GEN_0; // @[PRNG.scala 61:23]
  assign _T_1 = state_15 ^ state_13; // @[LFSR.scala 15:41]
  assign _T_2 = _T_1 ^ state_12; // @[LFSR.scala 15:41]
  assign _T_3 = _T_2 ^ state_10; // @[LFSR.scala 15:41]
  assign _GEN_0 = io_increment ? _T_3 : state_0; // @[PRNG.scala 61:23]
  assign io_out_0 = state_0; // @[PRNG.scala 69:10]
  assign io_out_1 = state_1; // @[PRNG.scala 69:10]
  assign io_out_2 = state_2; // @[PRNG.scala 69:10]
  assign io_out_3 = state_3; // @[PRNG.scala 69:10]
  assign io_out_4 = state_4; // @[PRNG.scala 69:10]
  assign io_out_5 = state_5; // @[PRNG.scala 69:10]
  assign io_out_6 = state_6; // @[PRNG.scala 69:10]
  assign io_out_7 = state_7; // @[PRNG.scala 69:10]
  assign io_out_8 = state_8; // @[PRNG.scala 69:10]
  assign io_out_9 = state_9; // @[PRNG.scala 69:10]
  assign io_out_10 = state_10; // @[PRNG.scala 69:10]
  assign io_out_11 = state_11; // @[PRNG.scala 69:10]
  assign io_out_12 = state_12; // @[PRNG.scala 69:10]
  assign io_out_13 = state_13; // @[PRNG.scala 69:10]
  assign io_out_14 = state_14; // @[PRNG.scala 69:10]
  assign io_out_15 = state_15; // @[PRNG.scala 69:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  state_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    state_0 <= reset | _GEN_0;
    if (reset) begin
      state_1 <= 1'h0;
    end else if (io_increment) begin
      state_1 <= state_0;
    end
    if (reset) begin
      state_2 <= 1'h0;
    end else if (io_increment) begin
      state_2 <= state_1;
    end
    if (reset) begin
      state_3 <= 1'h0;
    end else if (io_increment) begin
      state_3 <= state_2;
    end
    if (reset) begin
      state_4 <= 1'h0;
    end else if (io_increment) begin
      state_4 <= state_3;
    end
    if (reset) begin
      state_5 <= 1'h0;
    end else if (io_increment) begin
      state_5 <= state_4;
    end
    if (reset) begin
      state_6 <= 1'h0;
    end else if (io_increment) begin
      state_6 <= state_5;
    end
    if (reset) begin
      state_7 <= 1'h0;
    end else if (io_increment) begin
      state_7 <= state_6;
    end
    if (reset) begin
      state_8 <= 1'h0;
    end else if (io_increment) begin
      state_8 <= state_7;
    end
    if (reset) begin
      state_9 <= 1'h0;
    end else if (io_increment) begin
      state_9 <= state_8;
    end
    if (reset) begin
      state_10 <= 1'h0;
    end else if (io_increment) begin
      state_10 <= state_9;
    end
    if (reset) begin
      state_11 <= 1'h0;
    end else if (io_increment) begin
      state_11 <= state_10;
    end
    if (reset) begin
      state_12 <= 1'h0;
    end else if (io_increment) begin
      state_12 <= state_11;
    end
    if (reset) begin
      state_13 <= 1'h0;
    end else if (io_increment) begin
      state_13 <= state_12;
    end
    if (reset) begin
      state_14 <= 1'h0;
    end else if (io_increment) begin
      state_14 <= state_13;
    end
    if (reset) begin
      state_15 <= 1'h0;
    end else if (io_increment) begin
      state_15 <= state_14;
    end
  end
endmodule
module AXI4StreamBIST(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  input         auto_stream_out_ready,
  output        auto_stream_out_valid,
  output [31:0] auto_stream_out_bits_data,
  output        auto_stream_out_bits_last
);
  wire  MaxPeriodFibonacciLFSR_clock; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_reset; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_increment; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_0; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_1; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_2; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_3; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_4; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_5; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_6; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_7; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_8; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_9; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_10; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_11; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_12; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_13; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_14; // @[PRNG.scala 82:22]
  wire  MaxPeriodFibonacciLFSR_io_out_15; // @[PRNG.scala 82:22]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg  enable; // @[AXI4StreamBIST.scala 32:25]
  reg [31:0] _RAND_0;
  reg  terminate; // @[AXI4StreamBIST.scala 33:28]
  reg [31:0] _RAND_1;
  reg  cntrOrLFSR; // @[AXI4StreamBIST.scala 34:29]
  reg [31:0] _RAND_2;
  reg  upOrdown; // @[AXI4StreamBIST.scala 35:27]
  reg [31:0] _RAND_3;
  wire  bistOn; // @[AXI4StreamBIST.scala 37:25]
  wire  _T_1; // @[AXI4StreamBIST.scala 40:35]
  wire [7:0] _T_9; // @[PRNG.scala 86:17]
  wire [15:0] lfsr; // @[PRNG.scala 86:17]
  reg [7:0] cnt; // @[AXI4StreamBIST.scala 42:22]
  reg [31:0] _RAND_4;
  wire  cntEn; // @[AXI4StreamBIST.scala 43:24]
  wire  _T_17; // @[AXI4StreamBIST.scala 47:24]
  wire  _T_18; // @[AXI4StreamBIST.scala 47:17]
  wire [7:0] _T_20; // @[AXI4StreamBIST.scala 52:20]
  wire [7:0] _T_22; // @[AXI4StreamBIST.scala 55:20]
  wire  _T_23; // @[AXI4StreamBIST.scala 60:28]
  wire [15:0] _T_25; // @[AXI4StreamBIST.scala 61:25]
  wire  _T_27; // @[RegisterRouter.scala 40:39]
  wire  _T_28; // @[RegisterRouter.scala 40:26]
  wire  _T_29; // @[RegisterRouter.scala 42:29]
  wire  _T_72_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_36; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_224; // @[Cat.scala 29:58]
  wire [5:0] _T_76; // @[RegisterRouter.scala 59:16]
  wire  _T_82; // @[RegisterRouter.scala 59:16]
  wire  _T_30; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_39; // @[OneHot.scala 65:12]
  wire [1:0] _T_41; // @[Misc.scala 200:81]
  wire  _T_42; // @[Misc.scala 204:21]
  wire  _T_45; // @[Misc.scala 209:20]
  wire  _T_47; // @[Misc.scala 213:38]
  wire  _T_48; // @[Misc.scala 213:29]
  wire  _T_50; // @[Misc.scala 213:38]
  wire  _T_51; // @[Misc.scala 213:29]
  wire  _T_54; // @[Misc.scala 209:20]
  wire  _T_55; // @[Misc.scala 212:27]
  wire  _T_56; // @[Misc.scala 213:38]
  wire  _T_57; // @[Misc.scala 213:29]
  wire  _T_58; // @[Misc.scala 212:27]
  wire  _T_59; // @[Misc.scala 213:38]
  wire  _T_60; // @[Misc.scala 213:29]
  wire  _T_61; // @[Misc.scala 212:27]
  wire  _T_62; // @[Misc.scala 213:38]
  wire  _T_63; // @[Misc.scala 213:29]
  wire  _T_64; // @[Misc.scala 212:27]
  wire  _T_65; // @[Misc.scala 213:38]
  wire  _T_66; // @[Misc.scala 213:29]
  wire [3:0] _T_69; // @[Cat.scala 29:58]
  wire [3:0] _T_71; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_94; // @[Bitwise.scala 72:12]
  wire [7:0] _T_96; // @[Bitwise.scala 72:12]
  wire [7:0] _T_98; // @[Bitwise.scala 72:12]
  wire [7:0] _T_100; // @[Bitwise.scala 72:12]
  wire [31:0] _T_103; // @[Cat.scala 29:58]
  wire  _T_235; // @[RegisterRouter.scala 59:16]
  wire [3:0] _T_225; // @[OneHot.scala 58:35]
  wire  _T_262; // @[RegisterRouter.scala 59:16]
  wire  _T_274; // @[RegisterRouter.scala 59:16]
  wire  _T_275; // @[RegisterRouter.scala 59:16]
  wire  _T_129; // @[RegisterRouter.scala 59:16]
  wire  _T_269; // @[RegisterRouter.scala 59:16]
  wire  _T_270; // @[RegisterRouter.scala 59:16]
  wire  _T_152; // @[RegisterRouter.scala 59:16]
  wire  _T_279; // @[RegisterRouter.scala 59:16]
  wire  _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_175; // @[RegisterRouter.scala 59:16]
  wire  _T_264; // @[RegisterRouter.scala 59:16]
  wire  _T_265; // @[RegisterRouter.scala 59:16]
  wire  _T_198; // @[RegisterRouter.scala 59:16]
  wire  _GEN_24; // @[MuxLiteral.scala 48:10]
  wire  _GEN_25; // @[MuxLiteral.scala 48:10]
  wire  _GEN_26; // @[MuxLiteral.scala 48:10]
  wire  _GEN_28; // @[MuxLiteral.scala 48:10]
  wire  _GEN_29; // @[MuxLiteral.scala 48:10]
  wire  _GEN_30; // @[MuxLiteral.scala 48:10]
  wire  _T_349; // @[RegisterRouter.scala 59:16]
  wire  _T_350_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_350_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_353; // @[RegisterRouter.scala 65:29]
  MaxPeriodFibonacciLFSR MaxPeriodFibonacciLFSR ( // @[PRNG.scala 82:22]
    .clock(MaxPeriodFibonacciLFSR_clock),
    .reset(MaxPeriodFibonacciLFSR_reset),
    .io_increment(MaxPeriodFibonacciLFSR_io_increment),
    .io_out_0(MaxPeriodFibonacciLFSR_io_out_0),
    .io_out_1(MaxPeriodFibonacciLFSR_io_out_1),
    .io_out_2(MaxPeriodFibonacciLFSR_io_out_2),
    .io_out_3(MaxPeriodFibonacciLFSR_io_out_3),
    .io_out_4(MaxPeriodFibonacciLFSR_io_out_4),
    .io_out_5(MaxPeriodFibonacciLFSR_io_out_5),
    .io_out_6(MaxPeriodFibonacciLFSR_io_out_6),
    .io_out_7(MaxPeriodFibonacciLFSR_io_out_7),
    .io_out_8(MaxPeriodFibonacciLFSR_io_out_8),
    .io_out_9(MaxPeriodFibonacciLFSR_io_out_9),
    .io_out_10(MaxPeriodFibonacciLFSR_io_out_10),
    .io_out_11(MaxPeriodFibonacciLFSR_io_out_11),
    .io_out_12(MaxPeriodFibonacciLFSR_io_out_12),
    .io_out_13(MaxPeriodFibonacciLFSR_io_out_13),
    .io_out_14(MaxPeriodFibonacciLFSR_io_out_14),
    .io_out_15(MaxPeriodFibonacciLFSR_io_out_15)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign bistOn = enable & auto_stream_out_ready; // @[AXI4StreamBIST.scala 37:25]
  assign _T_1 = ~cntrOrLFSR; // @[AXI4StreamBIST.scala 40:35]
  assign _T_9 = {MaxPeriodFibonacciLFSR_io_out_7,MaxPeriodFibonacciLFSR_io_out_6,MaxPeriodFibonacciLFSR_io_out_5,MaxPeriodFibonacciLFSR_io_out_4,MaxPeriodFibonacciLFSR_io_out_3,MaxPeriodFibonacciLFSR_io_out_2,MaxPeriodFibonacciLFSR_io_out_1,MaxPeriodFibonacciLFSR_io_out_0}; // @[PRNG.scala 86:17]
  assign lfsr = {MaxPeriodFibonacciLFSR_io_out_15,MaxPeriodFibonacciLFSR_io_out_14,MaxPeriodFibonacciLFSR_io_out_13,MaxPeriodFibonacciLFSR_io_out_12,MaxPeriodFibonacciLFSR_io_out_11,MaxPeriodFibonacciLFSR_io_out_10,MaxPeriodFibonacciLFSR_io_out_9,MaxPeriodFibonacciLFSR_io_out_8,_T_9}; // @[PRNG.scala 86:17]
  assign cntEn = bistOn & cntrOrLFSR; // @[AXI4StreamBIST.scala 43:24]
  assign _T_17 = cnt == 8'hff; // @[AXI4StreamBIST.scala 47:24]
  assign _T_18 = cntEn & _T_17; // @[AXI4StreamBIST.scala 47:17]
  assign _T_20 = cnt + 8'h1; // @[AXI4StreamBIST.scala 52:20]
  assign _T_22 = cnt - 8'h1; // @[AXI4StreamBIST.scala 55:20]
  assign _T_23 = ~terminate; // @[AXI4StreamBIST.scala 60:28]
  assign _T_25 = cntrOrLFSR ? {{8'd0}, cnt} : lfsr; // @[AXI4StreamBIST.scala 61:25]
  assign _T_27 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_28 = auto_mem_in_ar_valid | _T_27; // @[RegisterRouter.scala 40:26]
  assign _T_29 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_72_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_36 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_224 = {_T_36[3],_T_36[2]}; // @[Cat.scala 29:58]
  assign _T_76 = _T_36[7:2] & 6'h3c; // @[RegisterRouter.scala 59:16]
  assign _T_82 = _T_76 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_30 = _T_72_ready & _T_29; // @[RegisterRouter.scala 42:26]
  assign _T_39 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_41 = _T_39 | 2'h1; // @[Misc.scala 200:81]
  assign _T_42 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_45 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_47 = _T_41[1] & _T_45; // @[Misc.scala 213:38]
  assign _T_48 = _T_42 | _T_47; // @[Misc.scala 213:29]
  assign _T_50 = _T_41[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_51 = _T_42 | _T_50; // @[Misc.scala 213:29]
  assign _T_54 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_55 = _T_45 & _T_54; // @[Misc.scala 212:27]
  assign _T_56 = _T_41[0] & _T_55; // @[Misc.scala 213:38]
  assign _T_57 = _T_48 | _T_56; // @[Misc.scala 213:29]
  assign _T_58 = _T_45 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_59 = _T_41[0] & _T_58; // @[Misc.scala 213:38]
  assign _T_60 = _T_48 | _T_59; // @[Misc.scala 213:29]
  assign _T_61 = auto_mem_in_ar_bits_addr[1] & _T_54; // @[Misc.scala 212:27]
  assign _T_62 = _T_41[0] & _T_61; // @[Misc.scala 213:38]
  assign _T_63 = _T_51 | _T_62; // @[Misc.scala 213:29]
  assign _T_64 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_65 = _T_41[0] & _T_64; // @[Misc.scala 213:38]
  assign _T_66 = _T_51 | _T_65; // @[Misc.scala 213:29]
  assign _T_69 = {_T_66,_T_63,_T_60,_T_57}; // @[Cat.scala 29:58]
  assign _T_71 = auto_mem_in_ar_valid ? _T_69 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_94 = _T_71[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_96 = _T_71[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_98 = _T_71[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_100 = _T_71[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_103 = {_T_100,_T_98,_T_96,_T_94}; // @[Cat.scala 29:58]
  assign _T_235 = _T_28 & _T_72_ready; // @[RegisterRouter.scala 59:16]
  assign _T_225 = 4'h1 << _T_224; // @[OneHot.scala 58:35]
  assign _T_262 = _T_235 & _T_29; // @[RegisterRouter.scala 59:16]
  assign _T_274 = _T_262 & _T_225[2]; // @[RegisterRouter.scala 59:16]
  assign _T_275 = _T_274 & _T_82; // @[RegisterRouter.scala 59:16]
  assign _T_129 = _T_275 & _T_103[0]; // @[RegisterRouter.scala 59:16]
  assign _T_269 = _T_262 & _T_225[1]; // @[RegisterRouter.scala 59:16]
  assign _T_270 = _T_269 & _T_82; // @[RegisterRouter.scala 59:16]
  assign _T_152 = _T_270 & _T_103[0]; // @[RegisterRouter.scala 59:16]
  assign _T_279 = _T_262 & _T_225[3]; // @[RegisterRouter.scala 59:16]
  assign _T_280 = _T_279 & _T_82; // @[RegisterRouter.scala 59:16]
  assign _T_175 = _T_280 & _T_103[0]; // @[RegisterRouter.scala 59:16]
  assign _T_264 = _T_262 & _T_225[0]; // @[RegisterRouter.scala 59:16]
  assign _T_265 = _T_264 & _T_82; // @[RegisterRouter.scala 59:16]
  assign _T_198 = _T_265 & _T_103[0]; // @[RegisterRouter.scala 59:16]
  assign _GEN_24 = 2'h1 == _T_224 ? _T_82 : _T_82; // @[MuxLiteral.scala 48:10]
  assign _GEN_25 = 2'h2 == _T_224 ? _T_82 : _GEN_24; // @[MuxLiteral.scala 48:10]
  assign _GEN_26 = 2'h3 == _T_224 ? _T_82 : _GEN_25; // @[MuxLiteral.scala 48:10]
  assign _GEN_28 = 2'h1 == _T_224 ? terminate : enable; // @[MuxLiteral.scala 48:10]
  assign _GEN_29 = 2'h2 == _T_224 ? cntrOrLFSR : _GEN_28; // @[MuxLiteral.scala 48:10]
  assign _GEN_30 = 2'h3 == _T_224 ? upOrdown : _GEN_29; // @[MuxLiteral.scala 48:10]
  assign _T_349 = _GEN_26 & _GEN_30; // @[RegisterRouter.scala 59:16]
  assign _T_350_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_350_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_353 = ~_T_350_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_30 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_30 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_350_valid & _T_353; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_350_valid & _T_350_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_out_valid = enable & _T_23; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_data = {{16'd0}, _T_25}; // @[LazyModule.scala 173:49]
  assign auto_stream_out_bits_last = terminate; // @[LazyModule.scala 173:49]
  assign MaxPeriodFibonacciLFSR_clock = clock;
  assign MaxPeriodFibonacciLFSR_reset = reset;
  assign MaxPeriodFibonacciLFSR_io_increment = bistOn & _T_1; // @[PRNG.scala 85:23]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_27; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{31'd0}, _T_349}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_350_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  terminate = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cntrOrLFSR = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  upOrdown = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cnt = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable <= 1'h0;
    end else if (_T_198) begin
      enable <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      terminate <= 1'h0;
    end else if (_T_152) begin
      terminate <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      cntrOrLFSR <= 1'h0;
    end else if (_T_129) begin
      cntrOrLFSR <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      upOrdown <= 1'h0;
    end else if (_T_175) begin
      upOrdown <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      cnt <= 8'h0;
    end else if (_T_18) begin
      cnt <= 8'h0;
    end else if (cntEn) begin
      if (upOrdown) begin
        cnt <= _T_20;
      end else begin
        cnt <= _T_22;
      end
    end
  end
endmodule
module AXI4Splitter_1(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_3_ready,
  output        auto_stream_out_3_valid,
  output [31:0] auto_stream_out_3_bits_data,
  output        auto_stream_out_3_bits_last,
  input         auto_stream_out_2_ready,
  output        auto_stream_out_2_valid,
  output [31:0] auto_stream_out_2_bits_data,
  output        auto_stream_out_2_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_6; // @[RegisterRouter.scala 40:39]
  wire  _T_7; // @[RegisterRouter.scala 40:26]
  wire  _T_8; // @[RegisterRouter.scala 42:29]
  wire  _T_51_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_15; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_57; // @[RegisterRouter.scala 59:16]
  wire  _T_9; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_18; // @[OneHot.scala 65:12]
  wire [1:0] _T_20; // @[Misc.scala 200:81]
  wire  _T_21; // @[Misc.scala 204:21]
  wire  _T_24; // @[Misc.scala 209:20]
  wire  _T_26; // @[Misc.scala 213:38]
  wire  _T_27; // @[Misc.scala 213:29]
  wire  _T_29; // @[Misc.scala 213:38]
  wire  _T_30; // @[Misc.scala 213:29]
  wire  _T_33; // @[Misc.scala 209:20]
  wire  _T_34; // @[Misc.scala 212:27]
  wire  _T_35; // @[Misc.scala 213:38]
  wire  _T_36; // @[Misc.scala 213:29]
  wire  _T_37; // @[Misc.scala 212:27]
  wire  _T_38; // @[Misc.scala 213:38]
  wire  _T_39; // @[Misc.scala 213:29]
  wire  _T_40; // @[Misc.scala 212:27]
  wire  _T_41; // @[Misc.scala 213:38]
  wire  _T_42; // @[Misc.scala 213:29]
  wire  _T_43; // @[Misc.scala 212:27]
  wire  _T_44; // @[Misc.scala 213:38]
  wire  _T_45; // @[Misc.scala 213:29]
  wire [3:0] _T_48; // @[Cat.scala 29:58]
  wire [3:0] _T_50; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [7:0] _T_75; // @[Bitwise.scala 72:12]
  wire [31:0] _T_78; // @[Cat.scala 29:58]
  wire  _T_97; // @[RegisterRouter.scala 59:16]
  wire  _T_150; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_144; // @[OneHot.scala 58:35]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_174; // @[RegisterRouter.scala 59:16]
  wire  _T_175; // @[RegisterRouter.scala 59:16]
  wire  _T_104; // @[RegisterRouter.scala 59:16]
  wire  _T_169; // @[RegisterRouter.scala 59:16]
  wire  _T_170; // @[RegisterRouter.scala 59:16]
  wire  _T_127; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_225_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_225_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_228; // @[RegisterRouter.scala 65:29]
  wire  _T_231; // @[Splitter.scala 45:34]
  wire  _T_232; // @[Splitter.scala 45:34]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  _T_233; // @[Splitter.scala 46:34]
  wire  _T_234; // @[Splitter.scala 46:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_235; // @[Splitter.scala 49:19]
  wire  _T_236; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_239; // @[Splitter.scala 62:34]
  wire  _T_243; // @[Splitter.scala 62:34]
  wire  _T_247; // @[Splitter.scala 62:34]
  wire  _T_251; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_6 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_7 = auto_mem_in_ar_valid | _T_6; // @[RegisterRouter.scala 40:26]
  assign _T_8 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_51_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_15 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_55 = _T_15[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_57 = _T_55 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_9 = _T_51_ready & _T_8; // @[RegisterRouter.scala 42:26]
  assign _T_18 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_20 = _T_18 | 2'h1; // @[Misc.scala 200:81]
  assign _T_21 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_24 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_26 = _T_20[1] & _T_24; // @[Misc.scala 213:38]
  assign _T_27 = _T_21 | _T_26; // @[Misc.scala 213:29]
  assign _T_29 = _T_20[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_30 = _T_21 | _T_29; // @[Misc.scala 213:29]
  assign _T_33 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_34 = _T_24 & _T_33; // @[Misc.scala 212:27]
  assign _T_35 = _T_20[0] & _T_34; // @[Misc.scala 213:38]
  assign _T_36 = _T_27 | _T_35; // @[Misc.scala 213:29]
  assign _T_37 = _T_24 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_38 = _T_20[0] & _T_37; // @[Misc.scala 213:38]
  assign _T_39 = _T_27 | _T_38; // @[Misc.scala 213:29]
  assign _T_40 = auto_mem_in_ar_bits_addr[1] & _T_33; // @[Misc.scala 212:27]
  assign _T_41 = _T_20[0] & _T_40; // @[Misc.scala 213:38]
  assign _T_42 = _T_30 | _T_41; // @[Misc.scala 213:29]
  assign _T_43 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_44 = _T_20[0] & _T_43; // @[Misc.scala 213:38]
  assign _T_45 = _T_30 | _T_44; // @[Misc.scala 213:29]
  assign _T_48 = {_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58]
  assign _T_50 = auto_mem_in_ar_valid ? _T_48 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_69 = _T_50[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_50[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_50[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_75 = _T_50[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_78 = {_T_75,_T_73,_T_71,_T_69}; // @[Cat.scala 29:58]
  assign _T_97 = _T_78 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_150 = _T_7 & _T_51_ready; // @[RegisterRouter.scala 59:16]
  assign _T_144 = 2'h1 << _T_15[2]; // @[OneHot.scala 58:35]
  assign _T_167 = _T_150 & _T_8; // @[RegisterRouter.scala 59:16]
  assign _T_174 = _T_167 & _T_144[1]; // @[RegisterRouter.scala 59:16]
  assign _T_175 = _T_174 & _T_57; // @[RegisterRouter.scala 59:16]
  assign _T_104 = _T_175 & _T_97; // @[RegisterRouter.scala 59:16]
  assign _T_169 = _T_167 & _T_144[0]; // @[RegisterRouter.scala 59:16]
  assign _T_170 = _T_169 & _T_57; // @[RegisterRouter.scala 59:16]
  assign _T_127 = _T_170 & _T_97; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_15[2] ? _T_57 : _T_57; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_15[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_225_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_225_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_228 = ~_T_225_bits_read; // @[RegisterRouter.scala 65:29]
  assign _T_231 = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign _T_232 = _T_231 | auto_stream_out_2_ready; // @[Splitter.scala 45:34]
  assign readyOR = _T_232 | auto_stream_out_3_ready; // @[Splitter.scala 45:34]
  assign _T_233 = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_234 = _T_233 & auto_stream_out_2_ready; // @[Splitter.scala 46:34]
  assign readyAND = _T_234 & auto_stream_out_3_ready; // @[Splitter.scala 46:34]
  assign _T_235 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_236 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_236 & readyOR; // @[Splitter.scala 52:33]
  assign _T_239 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_243 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign _T_247 = ~maskReg[2]; // @[Splitter.scala 62:34]
  assign _T_251 = ~maskReg[3]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_9 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_9 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_225_valid & _T_228; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_225_valid & _T_225_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_235 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_3_valid = auto_stream_in_valid & _T_251; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_3_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_valid = auto_stream_in_valid & _T_247; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_2_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_243; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_239; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_6; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_225_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_127) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_104) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module AXI4StreamMux_3(
  input         clock,
  input         reset,
  output        auto_register_in_aw_ready,
  input         auto_register_in_aw_valid,
  input         auto_register_in_aw_bits_id,
  input  [29:0] auto_register_in_aw_bits_addr,
  output        auto_register_in_w_ready,
  input         auto_register_in_w_valid,
  input  [31:0] auto_register_in_w_bits_data,
  input  [3:0]  auto_register_in_w_bits_strb,
  input         auto_register_in_b_ready,
  output        auto_register_in_b_valid,
  output        auto_register_in_b_bits_id,
  output        auto_register_in_ar_ready,
  input         auto_register_in_ar_valid,
  input         auto_register_in_ar_bits_id,
  input  [29:0] auto_register_in_ar_bits_addr,
  input  [2:0]  auto_register_in_ar_bits_size,
  input         auto_register_in_r_ready,
  output        auto_register_in_r_valid,
  output        auto_register_in_r_bits_id,
  output [31:0] auto_register_in_r_bits_data,
  output        auto_stream_in_5_ready,
  input         auto_stream_in_5_valid,
  input  [31:0] auto_stream_in_5_bits_data,
  input         auto_stream_in_5_bits_last,
  output        auto_stream_in_4_ready,
  input         auto_stream_in_4_valid,
  input  [31:0] auto_stream_in_4_bits_data,
  input         auto_stream_in_4_bits_last,
  output        auto_stream_in_3_ready,
  input         auto_stream_in_3_valid,
  input  [31:0] auto_stream_in_3_bits_data,
  input         auto_stream_in_3_bits_last,
  output        auto_stream_in_2_ready,
  input         auto_stream_in_2_valid,
  input  [31:0] auto_stream_in_2_bits_data,
  input         auto_stream_in_2_bits_last,
  output        auto_stream_in_1_ready,
  input         auto_stream_in_1_valid,
  input  [31:0] auto_stream_in_1_bits_data,
  input         auto_stream_in_1_bits_last,
  output        auto_stream_in_0_ready,
  input         auto_stream_in_0_valid,
  input  [31:0] auto_stream_in_0_bits_data,
  input         auto_stream_in_0_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [2:0] sels_0; // @[Mux.scala 32:23]
  reg [31:0] _RAND_0;
  reg [2:0] sels_1; // @[Mux.scala 32:23]
  reg [31:0] _RAND_1;
  reg [2:0] sels_2; // @[Mux.scala 32:23]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Mux.scala 45:28]
  wire  _GEN_7; // @[Mux.scala 45:41]
  wire  _GEN_8; // @[Mux.scala 45:41]
  wire  _T_4; // @[Mux.scala 45:28]
  wire  _GEN_12; // @[Mux.scala 45:41]
  wire [31:0] _GEN_15; // @[Mux.scala 45:41]
  wire  _GEN_16; // @[Mux.scala 45:41]
  wire  _GEN_17; // @[Mux.scala 45:41]
  wire  _T_5; // @[Mux.scala 45:28]
  wire  _GEN_21; // @[Mux.scala 45:41]
  wire [31:0] _GEN_24; // @[Mux.scala 45:41]
  wire  _GEN_25; // @[Mux.scala 45:41]
  wire  _GEN_26; // @[Mux.scala 45:41]
  wire  _T_6; // @[Mux.scala 45:28]
  wire  _GEN_30; // @[Mux.scala 45:41]
  wire [31:0] _GEN_33; // @[Mux.scala 45:41]
  wire  _GEN_34; // @[Mux.scala 45:41]
  wire  _GEN_35; // @[Mux.scala 45:41]
  wire  _T_7; // @[Mux.scala 45:28]
  wire  _GEN_39; // @[Mux.scala 45:41]
  wire [31:0] _GEN_42; // @[Mux.scala 45:41]
  wire  _GEN_43; // @[Mux.scala 45:41]
  wire  _GEN_44; // @[Mux.scala 45:41]
  wire  _T_8; // @[Mux.scala 45:28]
  wire  _GEN_53; // @[Mux.scala 45:41]
  wire  _T_9; // @[Mux.scala 40:46]
  wire [2:0] _T_11; // @[Mux.scala 41:29]
  wire  _T_12; // @[Mux.scala 45:28]
  wire  _GEN_61; // @[Mux.scala 45:41]
  wire  _GEN_62; // @[Mux.scala 45:41]
  wire  _T_13; // @[Mux.scala 45:28]
  wire  _GEN_66; // @[Mux.scala 45:41]
  wire [31:0] _GEN_69; // @[Mux.scala 45:41]
  wire  _GEN_70; // @[Mux.scala 45:41]
  wire  _GEN_71; // @[Mux.scala 45:41]
  wire  _T_14; // @[Mux.scala 45:28]
  wire  _GEN_75; // @[Mux.scala 45:41]
  wire [31:0] _GEN_78; // @[Mux.scala 45:41]
  wire  _GEN_79; // @[Mux.scala 45:41]
  wire  _GEN_80; // @[Mux.scala 45:41]
  wire  _T_15; // @[Mux.scala 45:28]
  wire  _GEN_84; // @[Mux.scala 45:41]
  wire [31:0] _GEN_87; // @[Mux.scala 45:41]
  wire  _GEN_88; // @[Mux.scala 45:41]
  wire  _GEN_89; // @[Mux.scala 45:41]
  wire  _T_16; // @[Mux.scala 45:28]
  wire  _GEN_93; // @[Mux.scala 45:41]
  wire [31:0] _GEN_96; // @[Mux.scala 45:41]
  wire  _GEN_97; // @[Mux.scala 45:41]
  wire  _GEN_98; // @[Mux.scala 45:41]
  wire  _T_17; // @[Mux.scala 45:28]
  wire  _GEN_107; // @[Mux.scala 45:41]
  wire  _T_18; // @[Mux.scala 40:46]
  wire  _T_19; // @[Mux.scala 40:46]
  wire  _T_21; // @[Mux.scala 40:75]
  wire [2:0] _T_22; // @[Mux.scala 41:29]
  wire  _T_23; // @[Mux.scala 45:28]
  wire  _T_24; // @[Mux.scala 45:28]
  wire  _T_25; // @[Mux.scala 45:28]
  wire  _T_26; // @[Mux.scala 45:28]
  wire  _T_27; // @[Mux.scala 45:28]
  wire  _T_28; // @[Mux.scala 45:28]
  wire  _T_30; // @[RegisterRouter.scala 40:39]
  wire  _T_31; // @[RegisterRouter.scala 40:26]
  wire  _T_32; // @[RegisterRouter.scala 42:29]
  wire  _T_75_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_39; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_194; // @[Cat.scala 29:58]
  wire  _T_33; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_42; // @[OneHot.scala 65:12]
  wire [1:0] _T_44; // @[Misc.scala 200:81]
  wire  _T_45; // @[Misc.scala 204:21]
  wire  _T_48; // @[Misc.scala 209:20]
  wire  _T_50; // @[Misc.scala 213:38]
  wire  _T_51; // @[Misc.scala 213:29]
  wire  _T_53; // @[Misc.scala 213:38]
  wire  _T_54; // @[Misc.scala 213:29]
  wire  _T_57; // @[Misc.scala 209:20]
  wire  _T_58; // @[Misc.scala 212:27]
  wire  _T_59; // @[Misc.scala 213:38]
  wire  _T_60; // @[Misc.scala 213:29]
  wire  _T_61; // @[Misc.scala 212:27]
  wire  _T_62; // @[Misc.scala 213:38]
  wire  _T_63; // @[Misc.scala 213:29]
  wire  _T_64; // @[Misc.scala 212:27]
  wire  _T_65; // @[Misc.scala 213:38]
  wire  _T_66; // @[Misc.scala 213:29]
  wire  _T_67; // @[Misc.scala 212:27]
  wire  _T_68; // @[Misc.scala 213:38]
  wire  _T_69; // @[Misc.scala 213:29]
  wire [3:0] _T_72; // @[Cat.scala 29:58]
  wire [3:0] _T_74; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_95; // @[Bitwise.scala 72:12]
  wire [7:0] _T_97; // @[Bitwise.scala 72:12]
  wire [7:0] _T_99; // @[Bitwise.scala 72:12]
  wire [7:0] _T_101; // @[Bitwise.scala 72:12]
  wire [31:0] _T_104; // @[Cat.scala 29:58]
  wire  _T_123; // @[RegisterRouter.scala 59:16]
  wire  _T_205; // @[RegisterRouter.scala 59:16]
  wire [3:0] _T_195; // @[OneHot.scala 58:35]
  wire  _T_232; // @[RegisterRouter.scala 59:16]
  wire  _T_244; // @[RegisterRouter.scala 59:16]
  wire  _T_130; // @[RegisterRouter.scala 59:16]
  wire  _T_239; // @[RegisterRouter.scala 59:16]
  wire  _T_153; // @[RegisterRouter.scala 59:16]
  wire  _T_234; // @[RegisterRouter.scala 59:16]
  wire  _T_176; // @[RegisterRouter.scala 59:16]
  wire [2:0] _GEN_186; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_187; // @[MuxLiteral.scala 48:10]
  wire [2:0] _GEN_188; // @[MuxLiteral.scala 48:10]
  wire  _T_320_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_320_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_323; // @[RegisterRouter.scala 65:29]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_3 = sels_0 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_7 = _T_3 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_8 = _T_3 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_4 = sels_0 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_12 = _T_4 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_15 = _T_4 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_16 = _T_4 ? auto_stream_in_1_valid : _GEN_7; // @[Mux.scala 45:41]
  assign _GEN_17 = _T_4 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_5 = sels_0 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_21 = _T_5 ? auto_stream_in_2_bits_last : _GEN_12; // @[Mux.scala 45:41]
  assign _GEN_24 = _T_5 ? auto_stream_in_2_bits_data : _GEN_15; // @[Mux.scala 45:41]
  assign _GEN_25 = _T_5 ? auto_stream_in_2_valid : _GEN_16; // @[Mux.scala 45:41]
  assign _GEN_26 = _T_5 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_6 = sels_0 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_30 = _T_6 ? auto_stream_in_3_bits_last : _GEN_21; // @[Mux.scala 45:41]
  assign _GEN_33 = _T_6 ? auto_stream_in_3_bits_data : _GEN_24; // @[Mux.scala 45:41]
  assign _GEN_34 = _T_6 ? auto_stream_in_3_valid : _GEN_25; // @[Mux.scala 45:41]
  assign _GEN_35 = _T_6 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_7 = sels_0 == 3'h4; // @[Mux.scala 45:28]
  assign _GEN_39 = _T_7 ? auto_stream_in_4_bits_last : _GEN_30; // @[Mux.scala 45:41]
  assign _GEN_42 = _T_7 ? auto_stream_in_4_bits_data : _GEN_33; // @[Mux.scala 45:41]
  assign _GEN_43 = _T_7 ? auto_stream_in_4_valid : _GEN_34; // @[Mux.scala 45:41]
  assign _GEN_44 = _T_7 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_8 = sels_0 == 3'h5; // @[Mux.scala 45:28]
  assign _GEN_53 = _T_8 & auto_stream_out_0_ready; // @[Mux.scala 45:41]
  assign _T_9 = sels_0 == sels_1; // @[Mux.scala 40:46]
  assign _T_11 = _T_9 ? 3'h6 : sels_1; // @[Mux.scala 41:29]
  assign _T_12 = _T_11 == 3'h0; // @[Mux.scala 45:28]
  assign _GEN_61 = _T_12 & auto_stream_in_0_valid; // @[Mux.scala 45:41]
  assign _GEN_62 = _T_12 ? auto_stream_out_1_ready : _GEN_8; // @[Mux.scala 45:41]
  assign _T_13 = _T_11 == 3'h1; // @[Mux.scala 45:28]
  assign _GEN_66 = _T_13 ? auto_stream_in_1_bits_last : auto_stream_in_0_bits_last; // @[Mux.scala 45:41]
  assign _GEN_69 = _T_13 ? auto_stream_in_1_bits_data : auto_stream_in_0_bits_data; // @[Mux.scala 45:41]
  assign _GEN_70 = _T_13 ? auto_stream_in_1_valid : _GEN_61; // @[Mux.scala 45:41]
  assign _GEN_71 = _T_13 ? auto_stream_out_1_ready : _GEN_17; // @[Mux.scala 45:41]
  assign _T_14 = _T_11 == 3'h2; // @[Mux.scala 45:28]
  assign _GEN_75 = _T_14 ? auto_stream_in_2_bits_last : _GEN_66; // @[Mux.scala 45:41]
  assign _GEN_78 = _T_14 ? auto_stream_in_2_bits_data : _GEN_69; // @[Mux.scala 45:41]
  assign _GEN_79 = _T_14 ? auto_stream_in_2_valid : _GEN_70; // @[Mux.scala 45:41]
  assign _GEN_80 = _T_14 ? auto_stream_out_1_ready : _GEN_26; // @[Mux.scala 45:41]
  assign _T_15 = _T_11 == 3'h3; // @[Mux.scala 45:28]
  assign _GEN_84 = _T_15 ? auto_stream_in_3_bits_last : _GEN_75; // @[Mux.scala 45:41]
  assign _GEN_87 = _T_15 ? auto_stream_in_3_bits_data : _GEN_78; // @[Mux.scala 45:41]
  assign _GEN_88 = _T_15 ? auto_stream_in_3_valid : _GEN_79; // @[Mux.scala 45:41]
  assign _GEN_89 = _T_15 ? auto_stream_out_1_ready : _GEN_35; // @[Mux.scala 45:41]
  assign _T_16 = _T_11 == 3'h4; // @[Mux.scala 45:28]
  assign _GEN_93 = _T_16 ? auto_stream_in_4_bits_last : _GEN_84; // @[Mux.scala 45:41]
  assign _GEN_96 = _T_16 ? auto_stream_in_4_bits_data : _GEN_87; // @[Mux.scala 45:41]
  assign _GEN_97 = _T_16 ? auto_stream_in_4_valid : _GEN_88; // @[Mux.scala 45:41]
  assign _GEN_98 = _T_16 ? auto_stream_out_1_ready : _GEN_44; // @[Mux.scala 45:41]
  assign _T_17 = _T_11 == 3'h5; // @[Mux.scala 45:28]
  assign _GEN_107 = _T_17 ? auto_stream_out_1_ready : _GEN_53; // @[Mux.scala 45:41]
  assign _T_18 = sels_0 == sels_2; // @[Mux.scala 40:46]
  assign _T_19 = sels_1 == sels_2; // @[Mux.scala 40:46]
  assign _T_21 = _T_18 | _T_19; // @[Mux.scala 40:75]
  assign _T_22 = _T_21 ? 3'h6 : sels_2; // @[Mux.scala 41:29]
  assign _T_23 = _T_22 == 3'h0; // @[Mux.scala 45:28]
  assign _T_24 = _T_22 == 3'h1; // @[Mux.scala 45:28]
  assign _T_25 = _T_22 == 3'h2; // @[Mux.scala 45:28]
  assign _T_26 = _T_22 == 3'h3; // @[Mux.scala 45:28]
  assign _T_27 = _T_22 == 3'h4; // @[Mux.scala 45:28]
  assign _T_28 = _T_22 == 3'h5; // @[Mux.scala 45:28]
  assign _T_30 = auto_register_in_aw_valid & auto_register_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_31 = auto_register_in_ar_valid | _T_30; // @[RegisterRouter.scala 40:26]
  assign _T_32 = ~auto_register_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_75_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_39 = auto_register_in_ar_valid ? auto_register_in_ar_bits_addr : auto_register_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_194 = {_T_39[3],_T_39[2]}; // @[Cat.scala 29:58]
  assign _T_33 = _T_75_ready & _T_32; // @[RegisterRouter.scala 42:26]
  assign _T_42 = 2'h1 << auto_register_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_44 = _T_42 | 2'h1; // @[Misc.scala 200:81]
  assign _T_45 = auto_register_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_48 = ~auto_register_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_50 = _T_44[1] & _T_48; // @[Misc.scala 213:38]
  assign _T_51 = _T_45 | _T_50; // @[Misc.scala 213:29]
  assign _T_53 = _T_44[1] & auto_register_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_54 = _T_45 | _T_53; // @[Misc.scala 213:29]
  assign _T_57 = ~auto_register_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_58 = _T_48 & _T_57; // @[Misc.scala 212:27]
  assign _T_59 = _T_44[0] & _T_58; // @[Misc.scala 213:38]
  assign _T_60 = _T_51 | _T_59; // @[Misc.scala 213:29]
  assign _T_61 = _T_48 & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_62 = _T_44[0] & _T_61; // @[Misc.scala 213:38]
  assign _T_63 = _T_51 | _T_62; // @[Misc.scala 213:29]
  assign _T_64 = auto_register_in_ar_bits_addr[1] & _T_57; // @[Misc.scala 212:27]
  assign _T_65 = _T_44[0] & _T_64; // @[Misc.scala 213:38]
  assign _T_66 = _T_54 | _T_65; // @[Misc.scala 213:29]
  assign _T_67 = auto_register_in_ar_bits_addr[1] & auto_register_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_68 = _T_44[0] & _T_67; // @[Misc.scala 213:38]
  assign _T_69 = _T_54 | _T_68; // @[Misc.scala 213:29]
  assign _T_72 = {_T_69,_T_66,_T_63,_T_60}; // @[Cat.scala 29:58]
  assign _T_74 = auto_register_in_ar_valid ? _T_72 : auto_register_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_95 = _T_74[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_97 = _T_74[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_99 = _T_74[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_101 = _T_74[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_104 = {_T_101,_T_99,_T_97,_T_95}; // @[Cat.scala 29:58]
  assign _T_123 = _T_104[2:0] == 3'h7; // @[RegisterRouter.scala 59:16]
  assign _T_205 = _T_31 & _T_75_ready; // @[RegisterRouter.scala 59:16]
  assign _T_195 = 4'h1 << _T_194; // @[OneHot.scala 58:35]
  assign _T_232 = _T_205 & _T_32; // @[RegisterRouter.scala 59:16]
  assign _T_244 = _T_232 & _T_195[2]; // @[RegisterRouter.scala 59:16]
  assign _T_130 = _T_244 & _T_123; // @[RegisterRouter.scala 59:16]
  assign _T_239 = _T_232 & _T_195[1]; // @[RegisterRouter.scala 59:16]
  assign _T_153 = _T_239 & _T_123; // @[RegisterRouter.scala 59:16]
  assign _T_234 = _T_232 & _T_195[0]; // @[RegisterRouter.scala 59:16]
  assign _T_176 = _T_234 & _T_123; // @[RegisterRouter.scala 59:16]
  assign _GEN_186 = 2'h1 == _T_194 ? sels_1 : sels_0; // @[MuxLiteral.scala 48:10]
  assign _GEN_187 = 2'h2 == _T_194 ? sels_2 : _GEN_186; // @[MuxLiteral.scala 48:10]
  assign _GEN_188 = 2'h3 == _T_194 ? 3'h0 : _GEN_187; // @[MuxLiteral.scala 48:10]
  assign _T_320_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_320_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_323 = ~_T_320_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_register_in_aw_ready = _T_33 & auto_register_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_w_ready = _T_33 & auto_register_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_valid = _T_320_valid & _T_323; // @[LazyModule.scala 173:31]
  assign auto_register_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_valid = _T_320_valid & _T_320_bits_read; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_register_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_5_ready = _T_28 | _GEN_107; // @[LazyModule.scala 173:31]
  assign auto_stream_in_4_ready = _T_27 | _GEN_98; // @[LazyModule.scala 173:31]
  assign auto_stream_in_3_ready = _T_26 | _GEN_89; // @[LazyModule.scala 173:31]
  assign auto_stream_in_2_ready = _T_25 | _GEN_80; // @[LazyModule.scala 173:31]
  assign auto_stream_in_1_ready = _T_24 | _GEN_71; // @[LazyModule.scala 173:31]
  assign auto_stream_in_0_ready = _T_23 | _GEN_62; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = _T_17 ? auto_stream_in_5_valid : _GEN_97; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = _T_17 ? auto_stream_in_5_bits_data : _GEN_96; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = _T_17 ? auto_stream_in_5_bits_last : _GEN_93; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = _T_8 ? auto_stream_in_5_valid : _GEN_43; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = _T_8 ? auto_stream_in_5_bits_data : _GEN_42; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = _T_8 ? auto_stream_in_5_bits_last : _GEN_39; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_register_in_ar_valid | _T_30; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_register_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = {{29'd0}, _GEN_188}; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_register_in_ar_valid ? auto_register_in_ar_bits_id : auto_register_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_320_bits_read ? auto_register_in_r_ready : auto_register_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sels_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sels_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sels_2 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      sels_0 <= 3'h6;
    end else if (_T_176) begin
      sels_0 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_1 <= 3'h6;
    end else if (_T_153) begin
      sels_1 <= auto_register_in_w_bits_data[2:0];
    end
    if (reset) begin
      sels_2 <= 3'h6;
    end else if (_T_130) begin
      sels_2 <= auto_register_in_w_bits_data[2:0];
    end
  end
endmodule
module AXI4Splitter_2(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_stream_in_ready,
  input         auto_stream_in_valid,
  input  [31:0] auto_stream_in_bits_data,
  input         auto_stream_in_bits_last,
  input         auto_stream_out_1_ready,
  output        auto_stream_out_1_valid,
  output [31:0] auto_stream_out_1_bits_data,
  output        auto_stream_out_1_bits_last,
  input         auto_stream_out_0_ready,
  output        auto_stream_out_0_valid,
  output [31:0] auto_stream_out_0_bits_data,
  output        auto_stream_out_0_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [31:0] ctrlReg; // @[Splitter.scala 27:26]
  reg [31:0] _RAND_0;
  reg [31:0] maskReg; // @[Splitter.scala 28:26]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[RegisterRouter.scala 40:39]
  wire  _T_5; // @[RegisterRouter.scala 40:26]
  wire  _T_6; // @[RegisterRouter.scala 42:29]
  wire  _T_49_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_13; // @[RegisterRouter.scala 48:19]
  wire [1:0] _T_53; // @[RegisterRouter.scala 59:16]
  wire  _T_55; // @[RegisterRouter.scala 59:16]
  wire  _T_7; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_16; // @[OneHot.scala 65:12]
  wire [1:0] _T_18; // @[Misc.scala 200:81]
  wire  _T_19; // @[Misc.scala 204:21]
  wire  _T_22; // @[Misc.scala 209:20]
  wire  _T_24; // @[Misc.scala 213:38]
  wire  _T_25; // @[Misc.scala 213:29]
  wire  _T_27; // @[Misc.scala 213:38]
  wire  _T_28; // @[Misc.scala 213:29]
  wire  _T_31; // @[Misc.scala 209:20]
  wire  _T_32; // @[Misc.scala 212:27]
  wire  _T_33; // @[Misc.scala 213:38]
  wire  _T_34; // @[Misc.scala 213:29]
  wire  _T_35; // @[Misc.scala 212:27]
  wire  _T_36; // @[Misc.scala 213:38]
  wire  _T_37; // @[Misc.scala 213:29]
  wire  _T_38; // @[Misc.scala 212:27]
  wire  _T_39; // @[Misc.scala 213:38]
  wire  _T_40; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 212:27]
  wire  _T_42; // @[Misc.scala 213:38]
  wire  _T_43; // @[Misc.scala 213:29]
  wire [3:0] _T_46; // @[Cat.scala 29:58]
  wire [3:0] _T_48; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_67; // @[Bitwise.scala 72:12]
  wire [7:0] _T_69; // @[Bitwise.scala 72:12]
  wire [7:0] _T_71; // @[Bitwise.scala 72:12]
  wire [7:0] _T_73; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76; // @[Cat.scala 29:58]
  wire  _T_95; // @[RegisterRouter.scala 59:16]
  wire  _T_148; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_142; // @[OneHot.scala 58:35]
  wire  _T_165; // @[RegisterRouter.scala 59:16]
  wire  _T_172; // @[RegisterRouter.scala 59:16]
  wire  _T_173; // @[RegisterRouter.scala 59:16]
  wire  _T_102; // @[RegisterRouter.scala 59:16]
  wire  _T_167; // @[RegisterRouter.scala 59:16]
  wire  _T_168; // @[RegisterRouter.scala 59:16]
  wire  _T_125; // @[RegisterRouter.scala 59:16]
  wire  _GEN_11; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_13; // @[MuxLiteral.scala 48:10]
  wire  _T_223_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_223_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_226; // @[RegisterRouter.scala 65:29]
  wire  readyOR; // @[Splitter.scala 45:34]
  wire  readyAND; // @[Splitter.scala 46:34]
  wire  _T_229; // @[Splitter.scala 49:19]
  wire  _T_230; // @[Splitter.scala 52:24]
  wire  _GEN_14; // @[Splitter.scala 52:33]
  wire  _T_233; // @[Splitter.scala 62:34]
  wire  _T_237; // @[Splitter.scala 62:34]
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign _T_4 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_5 = auto_mem_in_ar_valid | _T_4; // @[RegisterRouter.scala 40:26]
  assign _T_6 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_49_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_13 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_53 = _T_13[3:2] & 2'h2; // @[RegisterRouter.scala 59:16]
  assign _T_55 = _T_53 == 2'h0; // @[RegisterRouter.scala 59:16]
  assign _T_7 = _T_49_ready & _T_6; // @[RegisterRouter.scala 42:26]
  assign _T_16 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_18 = _T_16 | 2'h1; // @[Misc.scala 200:81]
  assign _T_19 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_22 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_24 = _T_18[1] & _T_22; // @[Misc.scala 213:38]
  assign _T_25 = _T_19 | _T_24; // @[Misc.scala 213:29]
  assign _T_27 = _T_18[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_28 = _T_19 | _T_27; // @[Misc.scala 213:29]
  assign _T_31 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_32 = _T_22 & _T_31; // @[Misc.scala 212:27]
  assign _T_33 = _T_18[0] & _T_32; // @[Misc.scala 213:38]
  assign _T_34 = _T_25 | _T_33; // @[Misc.scala 213:29]
  assign _T_35 = _T_22 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_36 = _T_18[0] & _T_35; // @[Misc.scala 213:38]
  assign _T_37 = _T_25 | _T_36; // @[Misc.scala 213:29]
  assign _T_38 = auto_mem_in_ar_bits_addr[1] & _T_31; // @[Misc.scala 212:27]
  assign _T_39 = _T_18[0] & _T_38; // @[Misc.scala 213:38]
  assign _T_40 = _T_28 | _T_39; // @[Misc.scala 213:29]
  assign _T_41 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_42 = _T_18[0] & _T_41; // @[Misc.scala 213:38]
  assign _T_43 = _T_28 | _T_42; // @[Misc.scala 213:29]
  assign _T_46 = {_T_43,_T_40,_T_37,_T_34}; // @[Cat.scala 29:58]
  assign _T_48 = auto_mem_in_ar_valid ? _T_46 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_67 = _T_48[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_69 = _T_48[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_71 = _T_48[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_73 = _T_48[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_76 = {_T_73,_T_71,_T_69,_T_67}; // @[Cat.scala 29:58]
  assign _T_95 = _T_76 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_148 = _T_5 & _T_49_ready; // @[RegisterRouter.scala 59:16]
  assign _T_142 = 2'h1 << _T_13[2]; // @[OneHot.scala 58:35]
  assign _T_165 = _T_148 & _T_6; // @[RegisterRouter.scala 59:16]
  assign _T_172 = _T_165 & _T_142[1]; // @[RegisterRouter.scala 59:16]
  assign _T_173 = _T_172 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_102 = _T_173 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _T_167 = _T_165 & _T_142[0]; // @[RegisterRouter.scala 59:16]
  assign _T_168 = _T_167 & _T_55; // @[RegisterRouter.scala 59:16]
  assign _T_125 = _T_168 & _T_95; // @[RegisterRouter.scala 59:16]
  assign _GEN_11 = _T_13[2] ? _T_55 : _T_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_13 = _T_13[2] ? maskReg : ctrlReg; // @[MuxLiteral.scala 48:10]
  assign _T_223_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_223_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_226 = ~_T_223_bits_read; // @[RegisterRouter.scala 65:29]
  assign readyOR = auto_stream_out_0_ready | auto_stream_out_1_ready; // @[Splitter.scala 45:34]
  assign readyAND = auto_stream_out_0_ready & auto_stream_out_1_ready; // @[Splitter.scala 46:34]
  assign _T_229 = ctrlReg == 32'h0; // @[Splitter.scala 49:19]
  assign _T_230 = ctrlReg == 32'h1; // @[Splitter.scala 52:24]
  assign _GEN_14 = _T_230 & readyOR; // @[Splitter.scala 52:33]
  assign _T_233 = ~maskReg[0]; // @[Splitter.scala 62:34]
  assign _T_237 = ~maskReg[1]; // @[Splitter.scala 62:34]
  assign auto_mem_in_aw_ready = _T_7 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_7 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_223_valid & _T_226; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_223_valid & _T_223_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_stream_in_ready = _T_229 ? readyAND : _GEN_14; // @[LazyModule.scala 173:31]
  assign auto_stream_out_1_valid = auto_stream_in_valid & _T_237; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_1_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_valid = auto_stream_in_valid & _T_233; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_data = auto_stream_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_stream_out_0_bits_last = auto_stream_in_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_4; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_11 ? _GEN_13 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_223_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ctrlReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maskReg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ctrlReg <= 32'h0;
    end else if (_T_125) begin
      ctrlReg <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      maskReg <= 32'h0;
    end else if (_T_102) begin
      maskReg <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module Queue_12(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_14_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:0]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_14_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_14_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_2;
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[Decoupled.scala 240:27]
  wire  _GEN_22; // @[Decoupled.scala 237:18]
  wire  _GEN_21; // @[Decoupled.scala 237:18]
  wire  _T_11; // @[Decoupled.scala 227:16]
  wire  _T_12; // @[Decoupled.scala 231:19]
  assign _T_data__T_14_addr = 1'h0;
  assign _T_data__T_14_data = _T_data[_T_data__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = 1'h0;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_last__T_14_addr = 1'h0;
  assign _T_last__T_14_data = _T_last[_T_last__T_14_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = 1'h0;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = _T_3 ? _GEN_13 : _T_6;
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_22 = _T_3 ? _GEN_13 : _T_6; // @[Decoupled.scala 237:18]
  assign _GEN_21 = _T_3 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_11 = _GEN_22 != _GEN_21; // @[Decoupled.scala 227:16]
  assign _T_12 = ~_T_3; // @[Decoupled.scala 231:19]
  assign io_enq_ready = io_deq_ready | _T_3; // @[Decoupled.scala 232:16 Decoupled.scala 245:40]
  assign io_deq_valid = io_enq_valid | _T_12; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits_data = _T_3 ? io_enq_bits_data : _T_data__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
  assign io_deq_bits_last = _T_3 ? io_enq_bits_last : _T_last__T_14_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_11) begin
      if (_T_3) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module StreamBuffer_1(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_12 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module AXI4StreamWidthAdapater_1_to_4(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [7:0]  auto_out_bits_data,
  output        auto_out_bits_last
);
  reg [1:0] _T_5; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_0;
  wire  _T_6; // @[AXI4StreamWidthAdapter.scala 159:14]
  wire  _T_7; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_8; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_9; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir0; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_11; // @[AXI4StreamWidthAdapter.scala 167:22]
  reg [31:0] _RAND_1;
  wire  _T_13; // @[AXI4StreamWidthAdapter.scala 168:38]
  wire [2:0] _T_14; // @[AXI4StreamWidthAdapter.scala 168:60]
  wire [2:0] _T_15; // @[AXI4StreamWidthAdapter.scala 168:33]
  wire [2:0] _GEN_1; // @[AXI4StreamWidthAdapter.scala 168:21]
  wire  ir1; // @[AXI4StreamWidthAdapter.scala 170:60]
  reg [1:0] _T_20; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_2;
  wire  _T_22; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_23; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_24; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_2; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir2; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_27; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_30; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_31; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_3; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir3; // @[AXI4StreamWidthAdapter.scala 163:34]
  reg [1:0] _T_34; // @[AXI4StreamWidthAdapter.scala 158:22]
  reg [31:0] _RAND_4;
  wire  _T_36; // @[AXI4StreamWidthAdapter.scala 159:38]
  wire [2:0] _T_37; // @[AXI4StreamWidthAdapter.scala 159:60]
  wire [2:0] _T_38; // @[AXI4StreamWidthAdapter.scala 159:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 159:21]
  wire  ir4; // @[AXI4StreamWidthAdapter.scala 163:34]
  wire  _T_56; // @[AXI4StreamWidthAdapter.scala 46:16]
  wire  _T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_59; // @[AXI4StreamWidthAdapter.scala 46:11]
  wire  _T_60; // @[AXI4StreamWidthAdapter.scala 47:16]
  wire  _T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_63; // @[AXI4StreamWidthAdapter.scala 47:11]
  wire  _T_64; // @[AXI4StreamWidthAdapter.scala 48:16]
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_67; // @[AXI4StreamWidthAdapter.scala 48:11]
  wire  _T_68; // @[AXI4StreamWidthAdapter.scala 49:16]
  wire  _T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire  _T_71; // @[AXI4StreamWidthAdapter.scala 49:11]
  wire [7:0] _GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  wire [7:0] _GEN_7; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign _T_6 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 159:14]
  assign _T_7 = _T_5 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_8 = _T_5 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_9 = _T_7 ? 3'h0 : _T_8; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_0 = _T_6 ? _T_9 : {{1'd0}, _T_5}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir0 = _T_7 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_13 = _T_11 == 2'h3; // @[AXI4StreamWidthAdapter.scala 168:38]
  assign _T_14 = _T_11 + 2'h1; // @[AXI4StreamWidthAdapter.scala 168:60]
  assign _T_15 = _T_13 ? 3'h0 : _T_14; // @[AXI4StreamWidthAdapter.scala 168:33]
  assign _GEN_1 = _T_6 ? _T_15 : {{1'd0}, _T_11}; // @[AXI4StreamWidthAdapter.scala 168:21]
  assign ir1 = _T_13 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 170:60]
  assign _T_22 = _T_20 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_23 = _T_20 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_24 = _T_22 ? 3'h0 : _T_23; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_2 = _T_6 ? _T_24 : {{1'd0}, _T_20}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir2 = _T_22 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_29 = _T_27 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_30 = _T_27 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_31 = _T_29 ? 3'h0 : _T_30; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_3 = _T_6 ? _T_31 : {{1'd0}, _T_27}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir3 = _T_29 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_36 = _T_34 == 2'h3; // @[AXI4StreamWidthAdapter.scala 159:38]
  assign _T_37 = _T_34 + 2'h1; // @[AXI4StreamWidthAdapter.scala 159:60]
  assign _T_38 = _T_36 ? 3'h0 : _T_37; // @[AXI4StreamWidthAdapter.scala 159:33]
  assign _GEN_4 = _T_6 ? _T_38 : {{1'd0}, _T_34}; // @[AXI4StreamWidthAdapter.scala 159:21]
  assign ir4 = _T_36 & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 163:34]
  assign _T_56 = ir0 == ir1; // @[AXI4StreamWidthAdapter.scala 46:16]
  assign _T_58 = _T_56 | reset; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign _T_59 = ~_T_58; // @[AXI4StreamWidthAdapter.scala 46:11]
  assign _T_60 = ir0 == ir2; // @[AXI4StreamWidthAdapter.scala 47:16]
  assign _T_62 = _T_60 | reset; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign _T_63 = ~_T_62; // @[AXI4StreamWidthAdapter.scala 47:11]
  assign _T_64 = ir0 == ir3; // @[AXI4StreamWidthAdapter.scala 48:16]
  assign _T_66 = _T_64 | reset; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign _T_67 = ~_T_66; // @[AXI4StreamWidthAdapter.scala 48:11]
  assign _T_68 = ir0 == ir4; // @[AXI4StreamWidthAdapter.scala 49:16]
  assign _T_70 = _T_68 | reset; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign _T_71 = ~_T_70; // @[AXI4StreamWidthAdapter.scala 49:11]
  assign _GEN_6 = 2'h1 == _T_5 ? auto_in_bits_data[15:8] : auto_in_bits_data[7:0]; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign _GEN_7 = 2'h2 == _T_5 ? auto_in_bits_data[23:16] : _GEN_6; // @[AXI4StreamWidthAdapter.scala 54:19]
  assign auto_in_ready = _T_7 & auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = 2'h3 == _T_5 ? auto_in_bits_data[31:24] : _GEN_7; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last & _T_13; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_11 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_20 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_27 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_34 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_5 <= 2'h0;
    end else begin
      _T_5 <= _GEN_0[1:0];
    end
    if (reset) begin
      _T_11 <= 2'h0;
    end else begin
      _T_11 <= _GEN_1[1:0];
    end
    if (reset) begin
      _T_20 <= 2'h0;
    end else begin
      _T_20 <= _GEN_2[1:0];
    end
    if (reset) begin
      _T_27 <= 2'h0;
    end else begin
      _T_27 <= _GEN_3[1:0];
    end
    if (reset) begin
      _T_34 <= 2'h0;
    end else begin
      _T_34 <= _GEN_4[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_59) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:46 assert(ir0 === ir1)\n"); // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_59) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 46:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:47 assert(ir0 === ir2)\n"); // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_63) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 47:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_67) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:48 assert(ir0 === ir3)\n"); // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_67) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 48:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_71) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:49 assert(ir0 === ir4)\n"); // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_71) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 49:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_13(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:3]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire [1:0] _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12; // @[Counter.scala 39:22]
  wire [1:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module StreamBuffer_2(
  input         clock,
  input         reset,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [31:0] auto_out_out_bits_data,
  output        auto_out_out_bits_last,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [31:0] auto_in_in_bits_data,
  input         auto_in_in_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_13 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_out_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign auto_in_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_out_ready; // @[Decoupled.scala 311:15]
endmodule
module AXI4StreamWidthAdapater_4_to_1_1(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [7:0]  auto_in_bits_data,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data
);
  reg [7:0] _T; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2; // @[AXI4StreamWidthAdapter.scala 101:37]
  reg [31:0] _RAND_2;
  reg [1:0] _T_3; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_3;
  wire  _T_4; // @[AXI4StreamWidthAdapter.scala 103:14]
  wire  _T_5; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_6; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_7; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_0; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  _T_9; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_10; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_12; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_13; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire  _T_15; // @[AXI4StreamWidthAdapter.scala 106:29]
  wire  _T_16; // @[AXI4StreamWidthAdapter.scala 106:22]
  wire [23:0] _T_18; // @[Cat.scala 29:58]
  wire  ov0; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_23; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_4;
  wire  _T_25; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_26; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_27; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_4; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov1; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_44; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_5;
  wire  _T_46; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_47; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_48; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_8; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov2; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_64; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_6;
  wire  _T_66; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_67; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_68; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_12; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov3; // @[AXI4StreamWidthAdapter.scala 112:32]
  reg [1:0] _T_84; // @[AXI4StreamWidthAdapter.scala 102:22]
  reg [31:0] _RAND_7;
  wire  _T_86; // @[AXI4StreamWidthAdapter.scala 103:38]
  wire [2:0] _T_87; // @[AXI4StreamWidthAdapter.scala 103:60]
  wire [2:0] _T_88; // @[AXI4StreamWidthAdapter.scala 103:33]
  wire [2:0] _GEN_16; // @[AXI4StreamWidthAdapter.scala 103:21]
  wire  ov4; // @[AXI4StreamWidthAdapter.scala 112:32]
  wire  _T_101; // @[AXI4StreamWidthAdapter.scala 42:16]
  wire  _T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_104; // @[AXI4StreamWidthAdapter.scala 42:11]
  wire  _T_105; // @[AXI4StreamWidthAdapter.scala 43:16]
  wire  _T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_108; // @[AXI4StreamWidthAdapter.scala 43:11]
  wire  _T_109; // @[AXI4StreamWidthAdapter.scala 44:16]
  wire  _T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_112; // @[AXI4StreamWidthAdapter.scala 44:11]
  wire  _T_113; // @[AXI4StreamWidthAdapter.scala 45:16]
  wire  _T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  wire  _T_116; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_4 = auto_in_valid & auto_out_ready; // @[AXI4StreamWidthAdapter.scala 103:14]
  assign _T_5 = _T_3 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_6 = _T_3 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_7 = _T_5 ? 3'h0 : _T_6; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_0 = _T_4 ? _T_7 : {{1'd0}, _T_3}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign _T_9 = _T_3 == 2'h0; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_10 = _T_4 & _T_9; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_12 = _T_3 == 2'h1; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_13 = _T_4 & _T_12; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_15 = _T_3 == 2'h2; // @[AXI4StreamWidthAdapter.scala 106:29]
  assign _T_16 = _T_4 & _T_15; // @[AXI4StreamWidthAdapter.scala 106:22]
  assign _T_18 = {auto_in_bits_data,_T_2,_T_1}; // @[Cat.scala 29:58]
  assign ov0 = _T_5 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_25 = _T_23 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_26 = _T_23 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_27 = _T_25 ? 3'h0 : _T_26; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_4 = _T_4 ? _T_27 : {{1'd0}, _T_23}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov1 = _T_25 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_46 = _T_44 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_47 = _T_44 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_48 = _T_46 ? 3'h0 : _T_47; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_8 = _T_4 ? _T_48 : {{1'd0}, _T_44}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov2 = _T_46 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_66 = _T_64 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_67 = _T_64 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_68 = _T_66 ? 3'h0 : _T_67; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_12 = _T_4 ? _T_68 : {{1'd0}, _T_64}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov3 = _T_66 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_86 = _T_84 == 2'h3; // @[AXI4StreamWidthAdapter.scala 103:38]
  assign _T_87 = _T_84 + 2'h1; // @[AXI4StreamWidthAdapter.scala 103:60]
  assign _T_88 = _T_86 ? 3'h0 : _T_87; // @[AXI4StreamWidthAdapter.scala 103:33]
  assign _GEN_16 = _T_4 ? _T_88 : {{1'd0}, _T_84}; // @[AXI4StreamWidthAdapter.scala 103:21]
  assign ov4 = _T_86 & auto_in_valid; // @[AXI4StreamWidthAdapter.scala 112:32]
  assign _T_101 = ov0 == ov1; // @[AXI4StreamWidthAdapter.scala 42:16]
  assign _T_103 = _T_101 | reset; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_104 = ~_T_103; // @[AXI4StreamWidthAdapter.scala 42:11]
  assign _T_105 = ov0 == ov2; // @[AXI4StreamWidthAdapter.scala 43:16]
  assign _T_107 = _T_105 | reset; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_108 = ~_T_107; // @[AXI4StreamWidthAdapter.scala 43:11]
  assign _T_109 = ov0 == ov3; // @[AXI4StreamWidthAdapter.scala 44:16]
  assign _T_111 = _T_109 | reset; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_112 = ~_T_111; // @[AXI4StreamWidthAdapter.scala 44:11]
  assign _T_113 = ov0 == ov4; // @[AXI4StreamWidthAdapter.scala 45:16]
  assign _T_115 = _T_113 | reset; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign _T_116 = ~_T_115; // @[AXI4StreamWidthAdapter.scala 45:11]
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = _T_5 & auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = {_T_18,_T}; // @[LazyModule.scala 173:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_23 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_44 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_64 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_84 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_10) begin
      _T <= auto_in_bits_data;
    end
    if (_T_13) begin
      _T_1 <= auto_in_bits_data;
    end
    if (_T_16) begin
      _T_2 <= auto_in_bits_data;
    end
    if (reset) begin
      _T_3 <= 2'h0;
    end else begin
      _T_3 <= _GEN_0[1:0];
    end
    if (reset) begin
      _T_23 <= 2'h0;
    end else begin
      _T_23 <= _GEN_4[1:0];
    end
    if (reset) begin
      _T_44 <= 2'h0;
    end else begin
      _T_44 <= _GEN_8[1:0];
    end
    if (reset) begin
      _T_64 <= 2'h0;
    end else begin
      _T_64 <= _GEN_12[1:0];
    end
    if (reset) begin
      _T_84 <= 2'h0;
    end else begin
      _T_84 <= _GEN_16[1:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_104) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:42 assert(ov0 === ov1)\n"); // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_104) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 42:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_108) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:43 assert(ov0 === ov2)\n"); // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_108) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 43:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_112) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:44 assert(ov0 === ov3)\n"); // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_112) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 44:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_116) begin
          $fwrite(32'h80000002,"Assertion failed\n    at AXI4StreamWidthAdapter.scala:45 assert(ov0 === ov4)\n"); // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_116) begin
          $fatal; // @[AXI4StreamWidthAdapter.scala 45:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module IntToBundleBridge(
  input   auto_in_0,
  output  auto_out_0
);
  assign auto_out_0 = auto_in_0; // @[LazyModule.scala 173:49]
endmodule
module UARTTx(
  input         clock,
  input         reset,
  input         io_en,
  output        io_in_ready,
  input         io_in_valid,
  input  [7:0]  io_in_bits,
  output        io_out,
  input  [15:0] io_div,
  input         io_nstop
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 44:11]
  reg [15:0] prescaler; // @[UARTTx.scala 21:22]
  reg [31:0] _RAND_0;
  wire  pulse; // @[UARTTx.scala 22:26]
  reg [3:0] counter; // @[UARTTx.scala 25:20]
  reg [31:0] _RAND_1;
  reg [8:0] shifter; // @[UARTTx.scala 26:20]
  reg [31:0] _RAND_2;
  reg  out; // @[UARTTx.scala 27:16]
  reg [31:0] _RAND_3;
  wire  plusarg_tx; // @[UARTTx.scala 30:90]
  wire  busy; // @[UARTTx.scala 32:23]
  wire  _T; // @[UARTTx.scala 33:27]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[UARTTx.scala 36:11]
  wire  _T_6; // @[UARTTx.scala 38:22]
  wire [9:0] _T_9; // @[Cat.scala 29:58]
  wire  _T_10; // @[UARTTx.scala 55:19]
  wire [3:0] _T_12; // @[Mux.scala 27:72]
  wire [3:0] _T_13; // @[Mux.scala 27:72]
  wire [3:0] _T_14; // @[Mux.scala 27:72]
  wire [3:0] _T_17; // @[UARTTx.scala 55:53]
  wire [9:0] _GEN_0; // @[UARTTx.scala 38:37]
  wire [15:0] _T_20; // @[UARTTx.scala 59:78]
  wire  _T_22; // @[UARTTx.scala 61:15]
  wire [3:0] _T_24; // @[UARTTx.scala 62:24]
  wire [8:0] _T_26; // @[Cat.scala 29:58]
  wire [9:0] _GEN_4; // @[UARTTx.scala 61:24]
  wire  _GEN_5; // @[UARTTx.scala 61:24]
  plusarg_reader #(.FORMAT("uart_tx=%d"), .DEFAULT(1), .WIDTH(32)) plusarg_reader ( // @[PlusArg.scala 44:11]
    .out(plusarg_reader_out)
  );
  assign pulse = prescaler == 16'h0; // @[UARTTx.scala 22:26]
  assign plusarg_tx = plusarg_reader_out != 32'h0; // @[UARTTx.scala 30:90]
  assign busy = counter != 4'h0; // @[UARTTx.scala 32:23]
  assign _T = ~busy; // @[UARTTx.scala 33:27]
  assign _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = ~reset; // @[UARTTx.scala 36:11]
  assign _T_6 = _T_2 & plusarg_tx; // @[UARTTx.scala 38:22]
  assign _T_9 = {1'h1,io_in_bits,1'h0}; // @[Cat.scala 29:58]
  assign _T_10 = ~io_nstop; // @[UARTTx.scala 55:19]
  assign _T_12 = _T_10 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  assign _T_13 = io_nstop ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  assign _T_14 = _T_12 | _T_13; // @[Mux.scala 27:72]
  assign _T_17 = _T_14 - 4'h0; // @[UARTTx.scala 55:53]
  assign _GEN_0 = _T_6 ? _T_9 : {{1'd0}, shifter}; // @[UARTTx.scala 38:37]
  assign _T_20 = prescaler - 16'h1; // @[UARTTx.scala 59:78]
  assign _T_22 = pulse & busy; // @[UARTTx.scala 61:15]
  assign _T_24 = counter - 4'h1; // @[UARTTx.scala 62:24]
  assign _T_26 = {1'h1,shifter[8:1]}; // @[Cat.scala 29:58]
  assign _GEN_4 = _T_22 ? {{1'd0}, _T_26} : _GEN_0; // @[UARTTx.scala 61:24]
  assign _GEN_5 = _T_22 ? shifter[0] : out; // @[UARTTx.scala 61:24]
  assign io_in_ready = io_en & _T; // @[UARTTx.scala 33:15]
  assign io_out = out; // @[UARTTx.scala 28:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prescaler = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  shifter = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      prescaler <= 16'h0;
    end else if (busy) begin
      if (pulse) begin
        prescaler <= io_div;
      end else begin
        prescaler <= _T_20;
      end
    end
    if (reset) begin
      counter <= 4'h0;
    end else if (_T_22) begin
      counter <= _T_24;
    end else if (_T_6) begin
      counter <= _T_17;
    end
    shifter <= _GEN_4[8:0];
    out <= reset | _GEN_5;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & _T_4) begin
          $fwrite(32'h80000002,"UART TX (%x): %c\n",io_in_bits,io_in_bits); // @[UARTTx.scala 36:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module QueueCompatibility(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  output [8:0] io_count
);
  reg [7:0] _T [0:255]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire [7:0] _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [7:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire [7:0] _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg [7:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg [7:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire [7:0] _T_12; // @[Counter.scala 39:22]
  wire [7:0] _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire [7:0] _T_20; // @[Decoupled.scala 248:40]
  wire  _T_21; // @[Decoupled.scala 250:32]
  wire [8:0] _T_22; // @[Decoupled.scala 250:20]
  wire [8:0] _GEN_8; // @[Decoupled.scala 250:62]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 8'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 8'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign _T_20 = value - value_1; // @[Decoupled.scala 248:40]
  assign _T_21 = _T_1 & _T_2; // @[Decoupled.scala 250:32]
  assign _T_22 = _T_21 ? 9'h100 : 9'h0; // @[Decoupled.scala 250:20]
  assign _GEN_8 = {{1'd0}, _T_20}; // @[Decoupled.scala 250:62]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits = _T__T_18_data; // @[Decoupled.scala 233:15]
  assign io_count = _T_22 | _GEN_8; // @[Decoupled.scala 250:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    _T[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 8'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 8'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module UARTRx(
  input         clock,
  input         reset,
  input         io_en,
  input         io_in,
  output        io_out_valid,
  output [7:0]  io_out_bits,
  input  [15:0] io_div
);
  reg [1:0] debounce; // @[UARTRx.scala 22:21]
  reg [31:0] _RAND_0;
  wire  debounce_max; // @[UARTRx.scala 23:32]
  wire  debounce_min; // @[UARTRx.scala 24:32]
  reg [12:0] prescaler; // @[UARTRx.scala 26:22]
  reg [31:0] _RAND_1;
  wire  pulse; // @[UARTRx.scala 28:26]
  reg [3:0] data_count; // @[UARTRx.scala 32:23]
  reg [31:0] _RAND_2;
  wire  data_last; // @[UARTRx.scala 33:31]
  reg [3:0] sample_count; // @[UARTRx.scala 35:25]
  reg [31:0] _RAND_3;
  wire  sample_mid; // @[UARTRx.scala 36:34]
  wire [7:0] _T_1; // @[Cat.scala 29:58]
  wire [7:0] countdown; // @[UARTRx.scala 38:49]
  wire [3:0] remainder; // @[UARTRx.scala 43:25]
  wire  extend; // @[UARTRx.scala 44:30]
  reg  state; // @[UARTRx.scala 59:18]
  reg [31:0] _RAND_4;
  wire  _T_14; // @[Conditional.scala 37:30]
  wire  _T_21; // @[UARTRx.scala 66:13]
  wire  _GEN_8; // @[UARTRx.scala 66:21]
  wire  start; // @[Conditional.scala 40:58]
  wire  restore; // @[UARTRx.scala 45:23]
  wire [12:0] prescaler_in; // @[UARTRx.scala 46:25]
  wire  _T_4; // @[UARTRx.scala 47:51]
  wire  _T_5; // @[UARTRx.scala 47:42]
  wire [12:0] _GEN_41; // @[UARTRx.scala 47:37]
  wire [12:0] prescaler_next; // @[UARTRx.scala 47:37]
  reg [2:0] sample; // @[UARTRx.scala 49:19]
  reg [31:0] _RAND_5;
  wire  _T_10; // @[Misc.scala 165:48]
  wire  _T_11; // @[Misc.scala 165:48]
  wire  _T_12; // @[Misc.scala 166:22]
  wire  _T_13; // @[Misc.scala 165:48]
  wire  voter; // @[Misc.scala 166:22]
  reg [7:0] shifter; // @[UARTRx.scala 51:20]
  reg [31:0] _RAND_6;
  reg  valid; // @[UARTRx.scala 53:18]
  reg [31:0] _RAND_7;
  wire  _T_16; // @[UARTRx.scala 63:13]
  wire  _T_17; // @[UARTRx.scala 63:26]
  wire  _T_18; // @[UARTRx.scala 63:23]
  wire [1:0] _T_20; // @[UARTRx.scala 64:30]
  wire [1:0] _T_23; // @[UARTRx.scala 67:30]
  wire [3:0] _T_27; // @[UARTRx.scala 72:94]
  wire  _GEN_1; // @[UARTRx.scala 68:29]
  wire [3:0] _T_29; // @[Cat.scala 29:58]
  wire [7:0] _T_33; // @[Cat.scala 29:58]
  wire  _GEN_16; // @[UARTRx.scala 85:27]
  wire [3:0] _GEN_18; // @[UARTRx.scala 80:20]
  wire  _GEN_22; // @[UARTRx.scala 80:20]
  wire [3:0] _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_29; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_37; // @[Conditional.scala 40:58]
  wire  _T_34; // @[UARTRx.scala 112:9]
  assign debounce_max = debounce == 2'h3; // @[UARTRx.scala 23:32]
  assign debounce_min = debounce == 2'h0; // @[UARTRx.scala 24:32]
  assign pulse = prescaler == 13'h0; // @[UARTRx.scala 28:26]
  assign data_last = data_count == 4'h0; // @[UARTRx.scala 33:31]
  assign sample_mid = sample_count == 4'h7; // @[UARTRx.scala 36:34]
  assign _T_1 = {data_count,sample_count}; // @[Cat.scala 29:58]
  assign countdown = _T_1 - 8'h1; // @[UARTRx.scala 38:49]
  assign remainder = io_div[3:0]; // @[UARTRx.scala 43:25]
  assign extend = sample_count < remainder; // @[UARTRx.scala 44:30]
  assign _T_14 = ~state; // @[Conditional.scala 37:30]
  assign _T_21 = ~io_in; // @[UARTRx.scala 66:13]
  assign _GEN_8 = _T_21 & debounce_max; // @[UARTRx.scala 66:21]
  assign start = _T_14 & _GEN_8; // @[Conditional.scala 40:58]
  assign restore = start | pulse; // @[UARTRx.scala 45:23]
  assign prescaler_in = restore ? {{1'd0}, io_div[15:4]} : prescaler; // @[UARTRx.scala 46:25]
  assign _T_4 = restore & extend; // @[UARTRx.scala 47:51]
  assign _T_5 = _T_4 ? 1'h0 : 1'h1; // @[UARTRx.scala 47:42]
  assign _GEN_41 = {{12'd0}, _T_5}; // @[UARTRx.scala 47:37]
  assign prescaler_next = prescaler_in - _GEN_41; // @[UARTRx.scala 47:37]
  assign _T_10 = sample[0] & sample[1]; // @[Misc.scala 165:48]
  assign _T_11 = sample[0] & sample[2]; // @[Misc.scala 165:48]
  assign _T_12 = _T_10 | _T_11; // @[Misc.scala 166:22]
  assign _T_13 = sample[1] & sample[2]; // @[Misc.scala 165:48]
  assign voter = _T_12 | _T_13; // @[Misc.scala 166:22]
  assign _T_16 = ~_T_21; // @[UARTRx.scala 63:13]
  assign _T_17 = ~debounce_min; // @[UARTRx.scala 63:26]
  assign _T_18 = _T_16 & _T_17; // @[UARTRx.scala 63:23]
  assign _T_20 = debounce - 2'h1; // @[UARTRx.scala 64:30]
  assign _T_23 = debounce + 2'h1; // @[UARTRx.scala 67:30]
  assign _T_27 = 4'h9 - 4'h0; // @[UARTRx.scala 72:94]
  assign _GEN_1 = debounce_max | state; // @[UARTRx.scala 68:29]
  assign _T_29 = {sample,io_in}; // @[Cat.scala 29:58]
  assign _T_33 = {voter,shifter[7:1]}; // @[Cat.scala 29:58]
  assign _GEN_16 = sample_mid & data_last; // @[UARTRx.scala 85:27]
  assign _GEN_18 = pulse ? _T_29 : {{1'd0}, sample}; // @[UARTRx.scala 80:20]
  assign _GEN_22 = pulse & _GEN_16; // @[UARTRx.scala 80:20]
  assign _GEN_25 = state ? _GEN_18 : {{1'd0}, sample}; // @[Conditional.scala 39:67]
  assign _GEN_29 = state & _GEN_22; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_14 ? {{1'd0}, sample} : _GEN_25; // @[Conditional.scala 40:58]
  assign _T_34 = ~io_en; // @[UARTRx.scala 112:9]
  assign io_out_valid = valid; // @[UARTRx.scala 55:16]
  assign io_out_bits = shifter; // @[UARTRx.scala 56:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  debounce = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  prescaler = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_count = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sample_count = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sample = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  shifter = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  valid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      debounce <= 2'h0;
    end else if (_T_34) begin
      debounce <= 2'h0;
    end else if (_T_14) begin
      if (_T_21) begin
        debounce <= _T_23;
      end else if (_T_18) begin
        debounce <= _T_20;
      end
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          prescaler <= prescaler_next;
        end
      end
    end else if (state) begin
      prescaler <= prescaler_next;
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          data_count <= _T_27;
        end
      end
    end else if (state) begin
      if (pulse) begin
        data_count <= countdown[7:4];
      end
    end
    if (_T_14) begin
      if (_T_21) begin
        if (debounce_max) begin
          sample_count <= 4'hf;
        end
      end
    end else if (state) begin
      if (pulse) begin
        sample_count <= countdown[3:0];
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_14) begin
      if (_T_21) begin
        state <= _GEN_1;
      end
    end else if (state) begin
      if (pulse) begin
        if (sample_mid) begin
          if (data_last) begin
            state <= 1'h0;
          end
        end
      end
    end
    sample <= _GEN_37[2:0];
    if (!(_T_14)) begin
      if (state) begin
        if (pulse) begin
          if (sample_mid) begin
            if (!(data_last)) begin
              shifter <= _T_33;
            end
          end
        end
      end
    end
    if (reset) begin
      valid <= 1'h0;
    end else if (_T_14) begin
      valid <= 1'h0;
    end else begin
      valid <= _GEN_29;
    end
  end
endmodule
module AXI4UARTBlock(
  input         clock,
  input         reset,
  output        auto_mem_in_aw_ready,
  input         auto_mem_in_aw_valid,
  input         auto_mem_in_aw_bits_id,
  input  [29:0] auto_mem_in_aw_bits_addr,
  output        auto_mem_in_w_ready,
  input         auto_mem_in_w_valid,
  input  [31:0] auto_mem_in_w_bits_data,
  input  [3:0]  auto_mem_in_w_bits_strb,
  input         auto_mem_in_b_ready,
  output        auto_mem_in_b_valid,
  output        auto_mem_in_b_bits_id,
  output        auto_mem_in_ar_ready,
  input         auto_mem_in_ar_valid,
  input         auto_mem_in_ar_bits_id,
  input  [29:0] auto_mem_in_ar_bits_addr,
  input  [2:0]  auto_mem_in_ar_bits_size,
  input         auto_mem_in_r_ready,
  output        auto_mem_in_r_valid,
  output        auto_mem_in_r_bits_id,
  output [31:0] auto_mem_in_r_bits_data,
  output        auto_in_in_ready,
  input         auto_in_in_valid,
  input  [7:0]  auto_in_in_bits_data,
  input         auto_out_out_ready,
  output        auto_out_out_valid,
  output [7:0]  auto_out_out_bits_data,
  output        int_0,
  output        io_txd,
  input         io_rxd
);
  wire  converter_auto_in_0; // @[Nodes.scala 31:31]
  wire  converter_auto_out_0; // @[Nodes.scala 31:31]
  wire  txm_clock; // @[DSPBlockUART.scala 101:21]
  wire  txm_reset; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_en; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_in_ready; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_in_valid; // @[DSPBlockUART.scala 101:21]
  wire [7:0] txm_io_in_bits; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_out; // @[DSPBlockUART.scala 101:21]
  wire [15:0] txm_io_div; // @[DSPBlockUART.scala 101:21]
  wire  txm_io_nstop; // @[DSPBlockUART.scala 101:21]
  wire  txq_clock; // @[DSPBlockUART.scala 102:21]
  wire  txq_reset; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_enq_ready; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_enq_valid; // @[DSPBlockUART.scala 102:21]
  wire [7:0] txq_io_enq_bits; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_deq_ready; // @[DSPBlockUART.scala 102:21]
  wire  txq_io_deq_valid; // @[DSPBlockUART.scala 102:21]
  wire [7:0] txq_io_deq_bits; // @[DSPBlockUART.scala 102:21]
  wire [8:0] txq_io_count; // @[DSPBlockUART.scala 102:21]
  wire  rxm_clock; // @[DSPBlockUART.scala 104:21]
  wire  rxm_reset; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_en; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_in; // @[DSPBlockUART.scala 104:21]
  wire  rxm_io_out_valid; // @[DSPBlockUART.scala 104:21]
  wire [7:0] rxm_io_out_bits; // @[DSPBlockUART.scala 104:21]
  wire [15:0] rxm_io_div; // @[DSPBlockUART.scala 104:21]
  wire  rxq_clock; // @[DSPBlockUART.scala 105:21]
  wire  rxq_reset; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_enq_ready; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_enq_valid; // @[DSPBlockUART.scala 105:21]
  wire [7:0] rxq_io_enq_bits; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_deq_ready; // @[DSPBlockUART.scala 105:21]
  wire  rxq_io_deq_valid; // @[DSPBlockUART.scala 105:21]
  wire [7:0] rxq_io_deq_bits; // @[DSPBlockUART.scala 105:21]
  wire [8:0] rxq_io_count; // @[DSPBlockUART.scala 105:21]
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_extra; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_read; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_extra; // @[Decoupled.scala 287:21]
  reg [15:0] div; // @[DSPBlockUART.scala 107:18]
  reg [31:0] _RAND_0;
  reg  txen; // @[DSPBlockUART.scala 113:19]
  reg [31:0] _RAND_1;
  reg  rxen; // @[DSPBlockUART.scala 114:19]
  reg [31:0] _RAND_2;
  reg [8:0] txwm; // @[DSPBlockUART.scala 121:19]
  reg [31:0] _RAND_3;
  reg [8:0] rxwm; // @[DSPBlockUART.scala 122:19]
  reg [31:0] _RAND_4;
  reg  nstop; // @[DSPBlockUART.scala 123:20]
  reg [31:0] _RAND_5;
  reg  ie_rxwm; // @[DSPBlockUART.scala 166:17]
  reg [31:0] _RAND_6;
  reg  ie_txwm; // @[DSPBlockUART.scala 166:17]
  reg [31:0] _RAND_7;
  wire  ip_txwm; // @[DSPBlockUART.scala 169:30]
  wire  ip_rxwm; // @[DSPBlockUART.scala 170:30]
  wire  _T_8; // @[DSPBlockUART.scala 171:31]
  wire  _T_9; // @[DSPBlockUART.scala 171:55]
  reg [31:0] _T_11; // @[DSPBlockUART.scala 175:53]
  reg [31:0] _RAND_8;
  reg [31:0] _T_12; // @[DSPBlockUART.scala 177:53]
  reg [31:0] _RAND_9;
  wire  _T_14; // @[RegisterRouter.scala 40:39]
  wire  _T_15; // @[RegisterRouter.scala 40:26]
  wire  _T_16; // @[RegisterRouter.scala 42:29]
  wire  _T_59_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  wire [29:0] _T_23; // @[RegisterRouter.scala 48:19]
  wire [2:0] _T_413; // @[Cat.scala 29:58]
  wire [5:0] _T_63; // @[RegisterRouter.scala 59:16]
  wire  _T_71; // @[RegisterRouter.scala 59:16]
  wire  _T_17; // @[RegisterRouter.scala 42:26]
  wire [1:0] _T_26; // @[OneHot.scala 65:12]
  wire [1:0] _T_28; // @[Misc.scala 200:81]
  wire  _T_29; // @[Misc.scala 204:21]
  wire  _T_32; // @[Misc.scala 209:20]
  wire  _T_34; // @[Misc.scala 213:38]
  wire  _T_35; // @[Misc.scala 213:29]
  wire  _T_37; // @[Misc.scala 213:38]
  wire  _T_38; // @[Misc.scala 213:29]
  wire  _T_41; // @[Misc.scala 209:20]
  wire  _T_42; // @[Misc.scala 212:27]
  wire  _T_43; // @[Misc.scala 213:38]
  wire  _T_44; // @[Misc.scala 213:29]
  wire  _T_45; // @[Misc.scala 212:27]
  wire  _T_46; // @[Misc.scala 213:38]
  wire  _T_47; // @[Misc.scala 213:29]
  wire  _T_48; // @[Misc.scala 212:27]
  wire  _T_49; // @[Misc.scala 213:38]
  wire  _T_50; // @[Misc.scala 213:29]
  wire  _T_51; // @[Misc.scala 212:27]
  wire  _T_52; // @[Misc.scala 213:38]
  wire  _T_53; // @[Misc.scala 213:29]
  wire [3:0] _T_56; // @[Cat.scala 29:58]
  wire [3:0] _T_58; // @[RegisterRouter.scala 54:25]
  wire [7:0] _T_87; // @[Bitwise.scala 72:12]
  wire [7:0] _T_89; // @[Bitwise.scala 72:12]
  wire [7:0] _T_91; // @[Bitwise.scala 72:12]
  wire [7:0] _T_93; // @[Bitwise.scala 72:12]
  wire [31:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_115; // @[RegisterRouter.scala 59:16]
  wire  _T_432; // @[RegisterRouter.scala 59:16]
  wire [7:0] _T_414; // @[OneHot.scala 58:35]
  wire  _T_479; // @[RegisterRouter.scala 59:16]
  wire  _T_481; // @[RegisterRouter.scala 59:16]
  wire  _T_482; // @[RegisterRouter.scala 59:16]
  wire  _T_122; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_180; // @[Cat.scala 29:58]
  wire  _T_486; // @[RegisterRouter.scala 59:16]
  wire  _T_487; // @[RegisterRouter.scala 59:16]
  wire  _T_193; // @[RegisterRouter.scala 59:16]
  wire  _T_209; // @[RegisterRouter.scala 59:16]
  wire  _T_511; // @[RegisterRouter.scala 59:16]
  wire  _T_512; // @[RegisterRouter.scala 59:16]
  wire  _T_216; // @[RegisterRouter.scala 59:16]
  wire  _T_491; // @[RegisterRouter.scala 59:16]
  wire  _T_492; // @[RegisterRouter.scala 59:16]
  wire  _T_239; // @[RegisterRouter.scala 59:16]
  wire  _T_262; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_274; // @[Cat.scala 29:58]
  wire  _T_280; // @[RegisterRouter.scala 59:16]
  wire  _T_287; // @[RegisterRouter.scala 59:16]
  wire [15:0] _T_298; // @[RegisterRouter.scala 59:16]
  wire [24:0] _T_299; // @[Cat.scala 29:58]
  wire  _T_496; // @[RegisterRouter.scala 59:16]
  wire  _T_497; // @[RegisterRouter.scala 59:16]
  wire  _T_312; // @[RegisterRouter.scala 59:16]
  wire  _T_335; // @[RegisterRouter.scala 59:16]
  wire [15:0] _T_346; // @[RegisterRouter.scala 59:16]
  wire [24:0] _T_347; // @[Cat.scala 29:58]
  wire  _T_501; // @[RegisterRouter.scala 59:16]
  wire  _T_502; // @[RegisterRouter.scala 59:16]
  wire  _T_360; // @[RegisterRouter.scala 59:16]
  wire  _T_383; // @[RegisterRouter.scala 59:16]
  wire [1:0] _T_395; // @[Cat.scala 29:58]
  wire  _GEN_43; // @[MuxLiteral.scala 48:10]
  wire  _GEN_44; // @[MuxLiteral.scala 48:10]
  wire  _GEN_45; // @[MuxLiteral.scala 48:10]
  wire  _GEN_46; // @[MuxLiteral.scala 48:10]
  wire  _GEN_47; // @[MuxLiteral.scala 48:10]
  wire  _GEN_48; // @[MuxLiteral.scala 48:10]
  wire  _GEN_58; // @[MuxLiteral.scala 48:10]
  wire  _GEN_49; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_51; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_2; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_52; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_3; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_53; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_4; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_54; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_5; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_55; // @[MuxLiteral.scala 48:10]
  wire [31:0] _T_624_6; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  wire [31:0] _GEN_56; // @[MuxLiteral.scala 48:10]
  wire [31:0] _GEN_57; // @[MuxLiteral.scala 48:10]
  wire  _T_627_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  wire  _T_627_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  wire  _T_630; // @[RegisterRouter.scala 65:29]
  IntToBundleBridge converter ( // @[Nodes.scala 31:31]
    .auto_in_0(converter_auto_in_0),
    .auto_out_0(converter_auto_out_0)
  );
  UARTTx txm ( // @[DSPBlockUART.scala 101:21]
    .clock(txm_clock),
    .reset(txm_reset),
    .io_en(txm_io_en),
    .io_in_ready(txm_io_in_ready),
    .io_in_valid(txm_io_in_valid),
    .io_in_bits(txm_io_in_bits),
    .io_out(txm_io_out),
    .io_div(txm_io_div),
    .io_nstop(txm_io_nstop)
  );
  QueueCompatibility txq ( // @[DSPBlockUART.scala 102:21]
    .clock(txq_clock),
    .reset(txq_reset),
    .io_enq_ready(txq_io_enq_ready),
    .io_enq_valid(txq_io_enq_valid),
    .io_enq_bits(txq_io_enq_bits),
    .io_deq_ready(txq_io_deq_ready),
    .io_deq_valid(txq_io_deq_valid),
    .io_deq_bits(txq_io_deq_bits),
    .io_count(txq_io_count)
  );
  UARTRx rxm ( // @[DSPBlockUART.scala 104:21]
    .clock(rxm_clock),
    .reset(rxm_reset),
    .io_en(rxm_io_en),
    .io_in(rxm_io_in),
    .io_out_valid(rxm_io_out_valid),
    .io_out_bits(rxm_io_out_bits),
    .io_div(rxm_io_div)
  );
  QueueCompatibility rxq ( // @[DSPBlockUART.scala 105:21]
    .clock(rxq_clock),
    .reset(rxq_reset),
    .io_enq_ready(rxq_io_enq_ready),
    .io_enq_valid(rxq_io_enq_valid),
    .io_enq_bits(rxq_io_enq_bits),
    .io_deq_ready(rxq_io_deq_ready),
    .io_deq_valid(rxq_io_deq_valid),
    .io_deq_bits(rxq_io_deq_bits),
    .io_count(rxq_io_count)
  );
  Queue Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign ip_txwm = txq_io_count < txwm; // @[DSPBlockUART.scala 169:30]
  assign ip_rxwm = rxq_io_count > rxwm; // @[DSPBlockUART.scala 170:30]
  assign _T_8 = ip_txwm & ie_txwm; // @[DSPBlockUART.scala 171:31]
  assign _T_9 = ip_rxwm & ie_rxwm; // @[DSPBlockUART.scala 171:55]
  assign _T_14 = auto_mem_in_aw_valid & auto_mem_in_w_valid; // @[RegisterRouter.scala 40:39]
  assign _T_15 = auto_mem_in_ar_valid | _T_14; // @[RegisterRouter.scala 40:26]
  assign _T_16 = ~auto_mem_in_ar_valid; // @[RegisterRouter.scala 42:29]
  assign _T_59_ready = Queue_io_enq_ready; // @[RegisterRouter.scala 59:16 Decoupled.scala 290:17]
  assign _T_23 = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_addr : auto_mem_in_aw_bits_addr; // @[RegisterRouter.scala 48:19]
  assign _T_413 = {_T_23[4],_T_23[3],_T_23[2]}; // @[Cat.scala 29:58]
  assign _T_63 = _T_23[7:2] & 6'h38; // @[RegisterRouter.scala 59:16]
  assign _T_71 = _T_63 == 6'h0; // @[RegisterRouter.scala 59:16]
  assign _T_17 = _T_59_ready & _T_16; // @[RegisterRouter.scala 42:26]
  assign _T_26 = 2'h1 << auto_mem_in_ar_bits_size[0]; // @[OneHot.scala 65:12]
  assign _T_28 = _T_26 | 2'h1; // @[Misc.scala 200:81]
  assign _T_29 = auto_mem_in_ar_bits_size >= 3'h2; // @[Misc.scala 204:21]
  assign _T_32 = ~auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 209:20]
  assign _T_34 = _T_28[1] & _T_32; // @[Misc.scala 213:38]
  assign _T_35 = _T_29 | _T_34; // @[Misc.scala 213:29]
  assign _T_37 = _T_28[1] & auto_mem_in_ar_bits_addr[1]; // @[Misc.scala 213:38]
  assign _T_38 = _T_29 | _T_37; // @[Misc.scala 213:29]
  assign _T_41 = ~auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 209:20]
  assign _T_42 = _T_32 & _T_41; // @[Misc.scala 212:27]
  assign _T_43 = _T_28[0] & _T_42; // @[Misc.scala 213:38]
  assign _T_44 = _T_35 | _T_43; // @[Misc.scala 213:29]
  assign _T_45 = _T_32 & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_46 = _T_28[0] & _T_45; // @[Misc.scala 213:38]
  assign _T_47 = _T_35 | _T_46; // @[Misc.scala 213:29]
  assign _T_48 = auto_mem_in_ar_bits_addr[1] & _T_41; // @[Misc.scala 212:27]
  assign _T_49 = _T_28[0] & _T_48; // @[Misc.scala 213:38]
  assign _T_50 = _T_38 | _T_49; // @[Misc.scala 213:29]
  assign _T_51 = auto_mem_in_ar_bits_addr[1] & auto_mem_in_ar_bits_addr[0]; // @[Misc.scala 212:27]
  assign _T_52 = _T_28[0] & _T_51; // @[Misc.scala 213:38]
  assign _T_53 = _T_38 | _T_52; // @[Misc.scala 213:29]
  assign _T_56 = {_T_53,_T_50,_T_47,_T_44}; // @[Cat.scala 29:58]
  assign _T_58 = auto_mem_in_ar_valid ? _T_56 : auto_mem_in_w_bits_strb; // @[RegisterRouter.scala 54:25]
  assign _T_87 = _T_58[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_89 = _T_58[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_91 = _T_58[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_93 = _T_58[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  assign _T_96 = {_T_93,_T_91,_T_89,_T_87}; // @[Cat.scala 29:58]
  assign _T_115 = _T_96 == 32'hffffffff; // @[RegisterRouter.scala 59:16]
  assign _T_432 = _T_15 & _T_59_ready; // @[RegisterRouter.scala 59:16]
  assign _T_414 = 8'h1 << _T_413; // @[OneHot.scala 58:35]
  assign _T_479 = _T_432 & _T_16; // @[RegisterRouter.scala 59:16]
  assign _T_481 = _T_479 & _T_414[0]; // @[RegisterRouter.scala 59:16]
  assign _T_482 = _T_481 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_122 = _T_482 & _T_115; // @[RegisterRouter.scala 59:16]
  assign _T_180 = {ip_rxwm,ip_txwm}; // @[Cat.scala 29:58]
  assign _T_486 = _T_479 & _T_414[1]; // @[RegisterRouter.scala 59:16]
  assign _T_487 = _T_486 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_193 = _T_487 & _T_115; // @[RegisterRouter.scala 59:16]
  assign _T_209 = _T_96[15:0] == 16'hffff; // @[RegisterRouter.scala 59:16]
  assign _T_511 = _T_479 & _T_414[6]; // @[RegisterRouter.scala 59:16]
  assign _T_512 = _T_511 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_216 = _T_512 & _T_209; // @[RegisterRouter.scala 59:16]
  assign _T_491 = _T_479 & _T_414[2]; // @[RegisterRouter.scala 59:16]
  assign _T_492 = _T_491 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_239 = _T_492 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  assign _T_262 = _T_492 & _T_96[1]; // @[RegisterRouter.scala 59:16]
  assign _T_274 = {nstop,txen}; // @[Cat.scala 29:58]
  assign _T_280 = _T_96[24:16] == 9'h1ff; // @[RegisterRouter.scala 59:16]
  assign _T_287 = _T_492 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_298 = {{14'd0}, _T_274}; // @[RegisterRouter.scala 59:16]
  assign _T_299 = {txwm,_T_298}; // @[Cat.scala 29:58]
  assign _T_496 = _T_479 & _T_414[3]; // @[RegisterRouter.scala 59:16]
  assign _T_497 = _T_496 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_312 = _T_497 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  assign _T_335 = _T_497 & _T_280; // @[RegisterRouter.scala 59:16]
  assign _T_346 = {{15'd0}, rxen}; // @[RegisterRouter.scala 59:16]
  assign _T_347 = {rxwm,_T_346}; // @[Cat.scala 29:58]
  assign _T_501 = _T_479 & _T_414[4]; // @[RegisterRouter.scala 59:16]
  assign _T_502 = _T_501 & _T_71; // @[RegisterRouter.scala 59:16]
  assign _T_360 = _T_502 & _T_96[0]; // @[RegisterRouter.scala 59:16]
  assign _T_383 = _T_502 & _T_96[1]; // @[RegisterRouter.scala 59:16]
  assign _T_395 = {ie_rxwm,ie_txwm}; // @[Cat.scala 29:58]
  assign _GEN_43 = 3'h1 == _T_413 ? _T_71 : _T_71; // @[MuxLiteral.scala 48:10]
  assign _GEN_44 = 3'h2 == _T_413 ? _T_71 : _GEN_43; // @[MuxLiteral.scala 48:10]
  assign _GEN_45 = 3'h3 == _T_413 ? _T_71 : _GEN_44; // @[MuxLiteral.scala 48:10]
  assign _GEN_46 = 3'h4 == _T_413 ? _T_71 : _GEN_45; // @[MuxLiteral.scala 48:10]
  assign _GEN_47 = 3'h5 == _T_413 ? _T_71 : _GEN_46; // @[MuxLiteral.scala 48:10]
  assign _GEN_48 = 3'h6 == _T_413 ? _T_71 : _GEN_47; // @[MuxLiteral.scala 48:10]
  assign _GEN_58 = 3'h7 == _T_413; // @[MuxLiteral.scala 48:10]
  assign _GEN_49 = _GEN_58 | _GEN_48; // @[MuxLiteral.scala 48:10]
  assign _GEN_51 = 3'h1 == _T_413 ? _T_12 : _T_11; // @[MuxLiteral.scala 48:10]
  assign _T_624_2 = {{7'd0}, _T_299}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_52 = 3'h2 == _T_413 ? _T_624_2 : _GEN_51; // @[MuxLiteral.scala 48:10]
  assign _T_624_3 = {{7'd0}, _T_347}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_53 = 3'h3 == _T_413 ? _T_624_3 : _GEN_52; // @[MuxLiteral.scala 48:10]
  assign _T_624_4 = {{30'd0}, _T_395}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_54 = 3'h4 == _T_413 ? _T_624_4 : _GEN_53; // @[MuxLiteral.scala 48:10]
  assign _T_624_5 = {{30'd0}, _T_180}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_55 = 3'h5 == _T_413 ? _T_624_5 : _GEN_54; // @[MuxLiteral.scala 48:10]
  assign _T_624_6 = {{16'd0}, div}; // @[MuxLiteral.scala 48:48 MuxLiteral.scala 48:48]
  assign _GEN_56 = 3'h6 == _T_413 ? _T_624_6 : _GEN_55; // @[MuxLiteral.scala 48:10]
  assign _GEN_57 = 3'h7 == _T_413 ? 32'h0 : _GEN_56; // @[MuxLiteral.scala 48:10]
  assign _T_627_bits_read = Queue_io_deq_bits_read; // @[Decoupled.scala 308:19 Decoupled.scala 309:14]
  assign _T_627_valid = Queue_io_deq_valid; // @[Decoupled.scala 308:19 Decoupled.scala 310:15]
  assign _T_630 = ~_T_627_bits_read; // @[RegisterRouter.scala 65:29]
  assign auto_mem_in_aw_ready = _T_17 & auto_mem_in_w_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_w_ready = _T_17 & auto_mem_in_aw_valid; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_valid = _T_627_valid & _T_630; // @[LazyModule.scala 173:31]
  assign auto_mem_in_b_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_ar_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_valid = _T_627_valid & _T_627_bits_read; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_id = Queue_io_deq_bits_extra; // @[LazyModule.scala 173:31]
  assign auto_mem_in_r_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_in_ready = txq_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_out_valid = rxq_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_out_bits_data = rxq_io_deq_bits; // @[LazyModule.scala 173:49]
  assign int_0 = converter_auto_out_0; // @[LISTestWithLA.scala 100:12]
  assign io_txd = txm_io_out; // @[DSPBlockUART.scala 135:12]
  assign converter_auto_in_0 = _T_8 | _T_9; // @[LazyModule.scala 167:57]
  assign txm_clock = clock;
  assign txm_reset = reset;
  assign txm_io_en = txen; // @[DSPBlockUART.scala 131:19]
  assign txm_io_in_valid = txq_io_deq_valid; // @[DSPBlockUART.scala 132:15]
  assign txm_io_in_bits = txq_io_deq_bits; // @[DSPBlockUART.scala 132:15]
  assign txm_io_div = div; // @[DSPBlockUART.scala 133:16]
  assign txm_io_nstop = nstop; // @[DSPBlockUART.scala 134:18]
  assign txq_clock = clock;
  assign txq_reset = reset;
  assign txq_io_enq_valid = auto_in_in_valid; // @[DSPBlockUART.scala 139:22]
  assign txq_io_enq_bits = auto_in_in_bits_data; // @[DSPBlockUART.scala 138:22]
  assign txq_io_deq_ready = txm_io_in_ready; // @[DSPBlockUART.scala 132:15]
  assign rxm_clock = clock;
  assign rxm_reset = reset;
  assign rxm_io_en = rxen; // @[DSPBlockUART.scala 151:15]
  assign rxm_io_in = io_rxd; // @[DSPBlockUART.scala 152:15]
  assign rxm_io_div = div; // @[DSPBlockUART.scala 154:16]
  assign rxq_clock = clock;
  assign rxq_reset = reset;
  assign rxq_io_enq_valid = rxm_io_out_valid; // @[DSPBlockUART.scala 153:16]
  assign rxq_io_enq_bits = rxm_io_out_bits; // @[DSPBlockUART.scala 153:16]
  assign rxq_io_deq_ready = auto_out_out_ready; // @[DSPBlockUART.scala 144:22]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_mem_in_ar_valid | _T_14; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_read = auto_mem_in_ar_valid; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_data = _GEN_49 ? _GEN_57 : 32'h0; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_extra = auto_mem_in_ar_valid ? auto_mem_in_ar_bits_id : auto_mem_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = _T_627_bits_read ? auto_mem_in_r_ready : auto_mem_in_b_ready; // @[Decoupled.scala 311:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  div = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  txen = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rxen = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  txwm = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rxwm = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  nstop = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ie_rxwm = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ie_txwm = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_11 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_12 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      div <= 16'had;
    end else if (_T_216) begin
      div <= auto_mem_in_w_bits_data[15:0];
    end
    if (reset) begin
      txen <= 1'h0;
    end else if (_T_239) begin
      txen <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      rxen <= 1'h0;
    end else if (_T_312) begin
      rxen <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      txwm <= 9'h0;
    end else if (_T_287) begin
      txwm <= auto_mem_in_w_bits_data[24:16];
    end
    if (reset) begin
      rxwm <= 9'h0;
    end else if (_T_335) begin
      rxwm <= auto_mem_in_w_bits_data[24:16];
    end
    if (reset) begin
      nstop <= 1'h0;
    end else if (_T_262) begin
      nstop <= auto_mem_in_w_bits_data[1];
    end
    if (reset) begin
      ie_rxwm <= 1'h0;
    end else if (_T_383) begin
      ie_rxwm <= auto_mem_in_w_bits_data[1];
    end
    if (reset) begin
      ie_txwm <= 1'h0;
    end else if (_T_360) begin
      ie_txwm <= auto_mem_in_w_bits_data[0];
    end
    if (reset) begin
      _T_11 <= 32'h0;
    end else if (_T_122) begin
      _T_11 <= auto_mem_in_w_bits_data;
    end
    if (reset) begin
      _T_12 <= 32'h0;
    end else if (_T_193) begin
      _T_12 <= auto_mem_in_w_bits_data;
    end
  end
endmodule
module QueueCompatibility_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [12:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [12:0] io_deq_bits
);
  reg [12:0] _T [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [12:0] _T__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T__T_18_addr; // @[Decoupled.scala 209:24]
  wire [12:0] _T__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_3;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _GEN_9; // @[Decoupled.scala 240:27]
  wire  _GEN_12; // @[Decoupled.scala 237:18]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _GEN_11; // @[Decoupled.scala 237:18]
  wire  _T_15; // @[Decoupled.scala 227:16]
  wire  _T_16; // @[Decoupled.scala 231:19]
  assign _T__T_18_addr = value_1;
  assign _T__T_18_data = _T[_T__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T__T_10_data = io_enq_bits;
  assign _T__T_10_addr = value;
  assign _T__T_10_mask = 1'h1;
  assign _T__T_10_en = _T_4 ? _GEN_9 : _T_6;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_6; // @[Decoupled.scala 240:27]
  assign _GEN_12 = _T_4 ? _GEN_9 : _T_6; // @[Decoupled.scala 237:18]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _GEN_11 = _T_4 ? 1'h0 : _T_8; // @[Decoupled.scala 237:18]
  assign _T_15 = _GEN_12 != _GEN_11; // @[Decoupled.scala 227:16]
  assign _T_16 = ~_T_4; // @[Decoupled.scala 231:19]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = io_enq_valid | _T_16; // @[Decoupled.scala 231:16 Decoupled.scala 236:40]
  assign io_deq_bits = _T_4 ? io_enq_bits : _T__T_18_data; // @[Decoupled.scala 233:15 Decoupled.scala 238:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T[initvar] = _RAND_0[12:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_10_en & _T__T_10_mask) begin
      _T[_T__T_10_addr] <= _T__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_GEN_12) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_GEN_11) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      if (_T_4) begin
        if (io_deq_ready) begin
          _T_1 <= 1'h0;
        end else begin
          _T_1 <= _T_6;
        end
      end else begin
        _T_1 <= _T_6;
      end
    end
  end
endmodule
module AXI4Xbar(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_12_aw_ready,
  output        auto_out_12_aw_valid,
  output        auto_out_12_aw_bits_id,
  output [29:0] auto_out_12_aw_bits_addr,
  output [2:0]  auto_out_12_aw_bits_size,
  input         auto_out_12_w_ready,
  output        auto_out_12_w_valid,
  output [31:0] auto_out_12_w_bits_data,
  output [3:0]  auto_out_12_w_bits_strb,
  output        auto_out_12_b_ready,
  input         auto_out_12_b_valid,
  input         auto_out_12_b_bits_id,
  input  [1:0]  auto_out_12_b_bits_resp,
  input         auto_out_12_ar_ready,
  output        auto_out_12_ar_valid,
  output        auto_out_12_ar_bits_id,
  output [29:0] auto_out_12_ar_bits_addr,
  output [2:0]  auto_out_12_ar_bits_size,
  output        auto_out_12_r_ready,
  input         auto_out_12_r_valid,
  input         auto_out_12_r_bits_id,
  input  [31:0] auto_out_12_r_bits_data,
  input  [1:0]  auto_out_12_r_bits_resp,
  input         auto_out_12_r_bits_last,
  input         auto_out_11_aw_ready,
  output        auto_out_11_aw_valid,
  output        auto_out_11_aw_bits_id,
  output [29:0] auto_out_11_aw_bits_addr,
  output [2:0]  auto_out_11_aw_bits_size,
  input         auto_out_11_w_ready,
  output        auto_out_11_w_valid,
  output [31:0] auto_out_11_w_bits_data,
  output [3:0]  auto_out_11_w_bits_strb,
  output        auto_out_11_b_ready,
  input         auto_out_11_b_valid,
  input         auto_out_11_b_bits_id,
  input  [1:0]  auto_out_11_b_bits_resp,
  input         auto_out_11_ar_ready,
  output        auto_out_11_ar_valid,
  output        auto_out_11_ar_bits_id,
  output [29:0] auto_out_11_ar_bits_addr,
  output [2:0]  auto_out_11_ar_bits_size,
  output        auto_out_11_r_ready,
  input         auto_out_11_r_valid,
  input         auto_out_11_r_bits_id,
  input  [31:0] auto_out_11_r_bits_data,
  input  [1:0]  auto_out_11_r_bits_resp,
  input         auto_out_11_r_bits_last,
  input         auto_out_10_aw_ready,
  output        auto_out_10_aw_valid,
  output        auto_out_10_aw_bits_id,
  output [29:0] auto_out_10_aw_bits_addr,
  output [2:0]  auto_out_10_aw_bits_size,
  input         auto_out_10_w_ready,
  output        auto_out_10_w_valid,
  output [31:0] auto_out_10_w_bits_data,
  output [3:0]  auto_out_10_w_bits_strb,
  output        auto_out_10_b_ready,
  input         auto_out_10_b_valid,
  input         auto_out_10_b_bits_id,
  input  [1:0]  auto_out_10_b_bits_resp,
  input         auto_out_10_ar_ready,
  output        auto_out_10_ar_valid,
  output        auto_out_10_ar_bits_id,
  output [29:0] auto_out_10_ar_bits_addr,
  output [2:0]  auto_out_10_ar_bits_size,
  output        auto_out_10_r_ready,
  input         auto_out_10_r_valid,
  input         auto_out_10_r_bits_id,
  input  [31:0] auto_out_10_r_bits_data,
  input  [1:0]  auto_out_10_r_bits_resp,
  input         auto_out_10_r_bits_last,
  input         auto_out_9_aw_ready,
  output        auto_out_9_aw_valid,
  output        auto_out_9_aw_bits_id,
  output [29:0] auto_out_9_aw_bits_addr,
  output [2:0]  auto_out_9_aw_bits_size,
  input         auto_out_9_w_ready,
  output        auto_out_9_w_valid,
  output [31:0] auto_out_9_w_bits_data,
  output [3:0]  auto_out_9_w_bits_strb,
  output        auto_out_9_b_ready,
  input         auto_out_9_b_valid,
  input         auto_out_9_b_bits_id,
  input  [1:0]  auto_out_9_b_bits_resp,
  input         auto_out_9_ar_ready,
  output        auto_out_9_ar_valid,
  output        auto_out_9_ar_bits_id,
  output [29:0] auto_out_9_ar_bits_addr,
  output [2:0]  auto_out_9_ar_bits_size,
  output        auto_out_9_r_ready,
  input         auto_out_9_r_valid,
  input         auto_out_9_r_bits_id,
  input  [31:0] auto_out_9_r_bits_data,
  input  [1:0]  auto_out_9_r_bits_resp,
  input         auto_out_9_r_bits_last,
  input         auto_out_8_aw_ready,
  output        auto_out_8_aw_valid,
  output        auto_out_8_aw_bits_id,
  output [29:0] auto_out_8_aw_bits_addr,
  output [2:0]  auto_out_8_aw_bits_size,
  input         auto_out_8_w_ready,
  output        auto_out_8_w_valid,
  output [31:0] auto_out_8_w_bits_data,
  output [3:0]  auto_out_8_w_bits_strb,
  output        auto_out_8_b_ready,
  input         auto_out_8_b_valid,
  input         auto_out_8_b_bits_id,
  input  [1:0]  auto_out_8_b_bits_resp,
  input         auto_out_8_ar_ready,
  output        auto_out_8_ar_valid,
  output        auto_out_8_ar_bits_id,
  output [29:0] auto_out_8_ar_bits_addr,
  output [2:0]  auto_out_8_ar_bits_size,
  output        auto_out_8_r_ready,
  input         auto_out_8_r_valid,
  input         auto_out_8_r_bits_id,
  input  [31:0] auto_out_8_r_bits_data,
  input  [1:0]  auto_out_8_r_bits_resp,
  input         auto_out_8_r_bits_last,
  input         auto_out_7_aw_ready,
  output        auto_out_7_aw_valid,
  output        auto_out_7_aw_bits_id,
  output [29:0] auto_out_7_aw_bits_addr,
  output [2:0]  auto_out_7_aw_bits_size,
  input         auto_out_7_w_ready,
  output        auto_out_7_w_valid,
  output [31:0] auto_out_7_w_bits_data,
  output [3:0]  auto_out_7_w_bits_strb,
  output        auto_out_7_b_ready,
  input         auto_out_7_b_valid,
  input         auto_out_7_b_bits_id,
  input  [1:0]  auto_out_7_b_bits_resp,
  input         auto_out_7_ar_ready,
  output        auto_out_7_ar_valid,
  output        auto_out_7_ar_bits_id,
  output [29:0] auto_out_7_ar_bits_addr,
  output [2:0]  auto_out_7_ar_bits_size,
  output        auto_out_7_r_ready,
  input         auto_out_7_r_valid,
  input         auto_out_7_r_bits_id,
  input  [31:0] auto_out_7_r_bits_data,
  input  [1:0]  auto_out_7_r_bits_resp,
  input         auto_out_7_r_bits_last,
  input         auto_out_6_aw_ready,
  output        auto_out_6_aw_valid,
  output        auto_out_6_aw_bits_id,
  output [29:0] auto_out_6_aw_bits_addr,
  output [2:0]  auto_out_6_aw_bits_size,
  input         auto_out_6_w_ready,
  output        auto_out_6_w_valid,
  output [31:0] auto_out_6_w_bits_data,
  output [3:0]  auto_out_6_w_bits_strb,
  output        auto_out_6_b_ready,
  input         auto_out_6_b_valid,
  input         auto_out_6_b_bits_id,
  input  [1:0]  auto_out_6_b_bits_resp,
  input         auto_out_6_ar_ready,
  output        auto_out_6_ar_valid,
  output        auto_out_6_ar_bits_id,
  output [29:0] auto_out_6_ar_bits_addr,
  output [2:0]  auto_out_6_ar_bits_size,
  output        auto_out_6_r_ready,
  input         auto_out_6_r_valid,
  input         auto_out_6_r_bits_id,
  input  [31:0] auto_out_6_r_bits_data,
  input  [1:0]  auto_out_6_r_bits_resp,
  input         auto_out_6_r_bits_last,
  input         auto_out_5_aw_ready,
  output        auto_out_5_aw_valid,
  output        auto_out_5_aw_bits_id,
  output [29:0] auto_out_5_aw_bits_addr,
  output [2:0]  auto_out_5_aw_bits_size,
  input         auto_out_5_w_ready,
  output        auto_out_5_w_valid,
  output [31:0] auto_out_5_w_bits_data,
  output [3:0]  auto_out_5_w_bits_strb,
  output        auto_out_5_b_ready,
  input         auto_out_5_b_valid,
  input         auto_out_5_b_bits_id,
  input  [1:0]  auto_out_5_b_bits_resp,
  input         auto_out_5_ar_ready,
  output        auto_out_5_ar_valid,
  output        auto_out_5_ar_bits_id,
  output [29:0] auto_out_5_ar_bits_addr,
  output [2:0]  auto_out_5_ar_bits_size,
  output        auto_out_5_r_ready,
  input         auto_out_5_r_valid,
  input         auto_out_5_r_bits_id,
  input  [31:0] auto_out_5_r_bits_data,
  input  [1:0]  auto_out_5_r_bits_resp,
  input         auto_out_5_r_bits_last,
  input         auto_out_4_aw_ready,
  output        auto_out_4_aw_valid,
  output        auto_out_4_aw_bits_id,
  output [29:0] auto_out_4_aw_bits_addr,
  output [2:0]  auto_out_4_aw_bits_size,
  input         auto_out_4_w_ready,
  output        auto_out_4_w_valid,
  output [31:0] auto_out_4_w_bits_data,
  output [3:0]  auto_out_4_w_bits_strb,
  output        auto_out_4_b_ready,
  input         auto_out_4_b_valid,
  input         auto_out_4_b_bits_id,
  input  [1:0]  auto_out_4_b_bits_resp,
  input         auto_out_4_ar_ready,
  output        auto_out_4_ar_valid,
  output        auto_out_4_ar_bits_id,
  output [29:0] auto_out_4_ar_bits_addr,
  output [2:0]  auto_out_4_ar_bits_size,
  output        auto_out_4_r_ready,
  input         auto_out_4_r_valid,
  input         auto_out_4_r_bits_id,
  input  [31:0] auto_out_4_r_bits_data,
  input  [1:0]  auto_out_4_r_bits_resp,
  input         auto_out_4_r_bits_last,
  input         auto_out_3_aw_ready,
  output        auto_out_3_aw_valid,
  output        auto_out_3_aw_bits_id,
  output [29:0] auto_out_3_aw_bits_addr,
  output [2:0]  auto_out_3_aw_bits_size,
  input         auto_out_3_w_ready,
  output        auto_out_3_w_valid,
  output [31:0] auto_out_3_w_bits_data,
  output [3:0]  auto_out_3_w_bits_strb,
  output        auto_out_3_b_ready,
  input         auto_out_3_b_valid,
  input         auto_out_3_b_bits_id,
  input  [1:0]  auto_out_3_b_bits_resp,
  input         auto_out_3_ar_ready,
  output        auto_out_3_ar_valid,
  output        auto_out_3_ar_bits_id,
  output [29:0] auto_out_3_ar_bits_addr,
  output [2:0]  auto_out_3_ar_bits_size,
  output        auto_out_3_r_ready,
  input         auto_out_3_r_valid,
  input         auto_out_3_r_bits_id,
  input  [31:0] auto_out_3_r_bits_data,
  input  [1:0]  auto_out_3_r_bits_resp,
  input         auto_out_3_r_bits_last,
  input         auto_out_2_aw_ready,
  output        auto_out_2_aw_valid,
  output        auto_out_2_aw_bits_id,
  output [29:0] auto_out_2_aw_bits_addr,
  output [2:0]  auto_out_2_aw_bits_size,
  input         auto_out_2_w_ready,
  output        auto_out_2_w_valid,
  output [31:0] auto_out_2_w_bits_data,
  output [3:0]  auto_out_2_w_bits_strb,
  output        auto_out_2_b_ready,
  input         auto_out_2_b_valid,
  input         auto_out_2_b_bits_id,
  input  [1:0]  auto_out_2_b_bits_resp,
  input         auto_out_2_ar_ready,
  output        auto_out_2_ar_valid,
  output        auto_out_2_ar_bits_id,
  output [29:0] auto_out_2_ar_bits_addr,
  output [2:0]  auto_out_2_ar_bits_size,
  output        auto_out_2_r_ready,
  input         auto_out_2_r_valid,
  input         auto_out_2_r_bits_id,
  input  [31:0] auto_out_2_r_bits_data,
  input  [1:0]  auto_out_2_r_bits_resp,
  input         auto_out_2_r_bits_last,
  input         auto_out_1_aw_ready,
  output        auto_out_1_aw_valid,
  output        auto_out_1_aw_bits_id,
  output [29:0] auto_out_1_aw_bits_addr,
  output [2:0]  auto_out_1_aw_bits_size,
  input         auto_out_1_w_ready,
  output        auto_out_1_w_valid,
  output [31:0] auto_out_1_w_bits_data,
  output [3:0]  auto_out_1_w_bits_strb,
  output        auto_out_1_b_ready,
  input         auto_out_1_b_valid,
  input         auto_out_1_b_bits_id,
  input  [1:0]  auto_out_1_b_bits_resp,
  input         auto_out_1_ar_ready,
  output        auto_out_1_ar_valid,
  output        auto_out_1_ar_bits_id,
  output [29:0] auto_out_1_ar_bits_addr,
  output [2:0]  auto_out_1_ar_bits_size,
  output        auto_out_1_r_ready,
  input         auto_out_1_r_valid,
  input         auto_out_1_r_bits_id,
  input  [31:0] auto_out_1_r_bits_data,
  input  [1:0]  auto_out_1_r_bits_resp,
  input         auto_out_1_r_bits_last,
  input         auto_out_0_aw_ready,
  output        auto_out_0_aw_valid,
  output        auto_out_0_aw_bits_id,
  output [29:0] auto_out_0_aw_bits_addr,
  output [2:0]  auto_out_0_aw_bits_size,
  input         auto_out_0_w_ready,
  output        auto_out_0_w_valid,
  output [31:0] auto_out_0_w_bits_data,
  output [3:0]  auto_out_0_w_bits_strb,
  output        auto_out_0_b_ready,
  input         auto_out_0_b_valid,
  input         auto_out_0_b_bits_id,
  input  [1:0]  auto_out_0_b_bits_resp,
  input         auto_out_0_ar_ready,
  output        auto_out_0_ar_valid,
  output        auto_out_0_ar_bits_id,
  output [29:0] auto_out_0_ar_bits_addr,
  output [2:0]  auto_out_0_ar_bits_size,
  output        auto_out_0_r_ready,
  input         auto_out_0_r_valid,
  input         auto_out_0_r_bits_id,
  input  [31:0] auto_out_0_r_bits_data,
  input  [1:0]  auto_out_0_r_bits_resp,
  input         auto_out_0_r_bits_last
);
  wire  awIn_0_clock; // @[Xbar.scala 55:47]
  wire  awIn_0_reset; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_enq_valid; // @[Xbar.scala 55:47]
  wire [12:0] awIn_0_io_enq_bits; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_ready; // @[Xbar.scala 55:47]
  wire  awIn_0_io_deq_valid; // @[Xbar.scala 55:47]
  wire [12:0] awIn_0_io_deq_bits; // @[Xbar.scala 55:47]
  wire [30:0] _T_1; // @[Parameters.scala 137:49]
  wire [30:0] _T_3; // @[Parameters.scala 137:52]
  wire  requestARIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_5; // @[Parameters.scala 137:31]
  wire [30:0] _T_6; // @[Parameters.scala 137:49]
  wire [30:0] _T_8; // @[Parameters.scala 137:52]
  wire  requestARIO_0_1; // @[Parameters.scala 137:67]
  wire [29:0] _T_10; // @[Parameters.scala 137:31]
  wire [30:0] _T_11; // @[Parameters.scala 137:49]
  wire [30:0] _T_13; // @[Parameters.scala 137:52]
  wire  requestARIO_0_2; // @[Parameters.scala 137:67]
  wire [29:0] _T_15; // @[Parameters.scala 137:31]
  wire [30:0] _T_16; // @[Parameters.scala 137:49]
  wire [30:0] _T_18; // @[Parameters.scala 137:52]
  wire  requestARIO_0_3; // @[Parameters.scala 137:67]
  wire [29:0] _T_20; // @[Parameters.scala 137:31]
  wire [30:0] _T_21; // @[Parameters.scala 137:49]
  wire [30:0] _T_23; // @[Parameters.scala 137:52]
  wire  requestARIO_0_4; // @[Parameters.scala 137:67]
  wire [29:0] _T_25; // @[Parameters.scala 137:31]
  wire [30:0] _T_26; // @[Parameters.scala 137:49]
  wire [30:0] _T_28; // @[Parameters.scala 137:52]
  wire  requestARIO_0_5; // @[Parameters.scala 137:67]
  wire [29:0] _T_30; // @[Parameters.scala 137:31]
  wire [30:0] _T_31; // @[Parameters.scala 137:49]
  wire [30:0] _T_33; // @[Parameters.scala 137:52]
  wire  requestARIO_0_6; // @[Parameters.scala 137:67]
  wire [29:0] _T_35; // @[Parameters.scala 137:31]
  wire [30:0] _T_36; // @[Parameters.scala 137:49]
  wire [30:0] _T_38; // @[Parameters.scala 137:52]
  wire  requestARIO_0_7; // @[Parameters.scala 137:67]
  wire [29:0] _T_40; // @[Parameters.scala 137:31]
  wire [30:0] _T_41; // @[Parameters.scala 137:49]
  wire [30:0] _T_43; // @[Parameters.scala 137:52]
  wire  requestARIO_0_8; // @[Parameters.scala 137:67]
  wire [29:0] _T_45; // @[Parameters.scala 137:31]
  wire [30:0] _T_46; // @[Parameters.scala 137:49]
  wire [30:0] _T_48; // @[Parameters.scala 137:52]
  wire  requestARIO_0_9; // @[Parameters.scala 137:67]
  wire [29:0] _T_50; // @[Parameters.scala 137:31]
  wire [30:0] _T_51; // @[Parameters.scala 137:49]
  wire [30:0] _T_53; // @[Parameters.scala 137:52]
  wire  requestARIO_0_10; // @[Parameters.scala 137:67]
  wire [29:0] _T_55; // @[Parameters.scala 137:31]
  wire [30:0] _T_56; // @[Parameters.scala 137:49]
  wire [30:0] _T_58; // @[Parameters.scala 137:52]
  wire  requestARIO_0_11; // @[Parameters.scala 137:67]
  wire [29:0] _T_60; // @[Parameters.scala 137:31]
  wire [30:0] _T_61; // @[Parameters.scala 137:49]
  wire [30:0] _T_63; // @[Parameters.scala 137:52]
  wire  requestARIO_0_12; // @[Parameters.scala 137:67]
  wire [30:0] _T_66; // @[Parameters.scala 137:49]
  wire [30:0] _T_68; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_0; // @[Parameters.scala 137:67]
  wire [29:0] _T_70; // @[Parameters.scala 137:31]
  wire [30:0] _T_71; // @[Parameters.scala 137:49]
  wire [30:0] _T_73; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_1; // @[Parameters.scala 137:67]
  wire [29:0] _T_75; // @[Parameters.scala 137:31]
  wire [30:0] _T_76; // @[Parameters.scala 137:49]
  wire [30:0] _T_78; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_2; // @[Parameters.scala 137:67]
  wire [29:0] _T_80; // @[Parameters.scala 137:31]
  wire [30:0] _T_81; // @[Parameters.scala 137:49]
  wire [30:0] _T_83; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_3; // @[Parameters.scala 137:67]
  wire [29:0] _T_85; // @[Parameters.scala 137:31]
  wire [30:0] _T_86; // @[Parameters.scala 137:49]
  wire [30:0] _T_88; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_4; // @[Parameters.scala 137:67]
  wire [29:0] _T_90; // @[Parameters.scala 137:31]
  wire [30:0] _T_91; // @[Parameters.scala 137:49]
  wire [30:0] _T_93; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_5; // @[Parameters.scala 137:67]
  wire [29:0] _T_95; // @[Parameters.scala 137:31]
  wire [30:0] _T_96; // @[Parameters.scala 137:49]
  wire [30:0] _T_98; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_6; // @[Parameters.scala 137:67]
  wire [29:0] _T_100; // @[Parameters.scala 137:31]
  wire [30:0] _T_101; // @[Parameters.scala 137:49]
  wire [30:0] _T_103; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_7; // @[Parameters.scala 137:67]
  wire [29:0] _T_105; // @[Parameters.scala 137:31]
  wire [30:0] _T_106; // @[Parameters.scala 137:49]
  wire [30:0] _T_108; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_8; // @[Parameters.scala 137:67]
  wire [29:0] _T_110; // @[Parameters.scala 137:31]
  wire [30:0] _T_111; // @[Parameters.scala 137:49]
  wire [30:0] _T_113; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_9; // @[Parameters.scala 137:67]
  wire [29:0] _T_115; // @[Parameters.scala 137:31]
  wire [30:0] _T_116; // @[Parameters.scala 137:49]
  wire [30:0] _T_118; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_10; // @[Parameters.scala 137:67]
  wire [29:0] _T_120; // @[Parameters.scala 137:31]
  wire [30:0] _T_121; // @[Parameters.scala 137:49]
  wire [30:0] _T_123; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_11; // @[Parameters.scala 137:67]
  wire [29:0] _T_125; // @[Parameters.scala 137:31]
  wire [30:0] _T_126; // @[Parameters.scala 137:49]
  wire [30:0] _T_128; // @[Parameters.scala 137:52]
  wire  requestAWIO_0_12; // @[Parameters.scala 137:67]
  wire  requestROI_0_0; // @[Parameters.scala 47:9]
  wire  requestROI_1_0; // @[Parameters.scala 47:9]
  wire  requestROI_2_0; // @[Parameters.scala 47:9]
  wire  requestROI_3_0; // @[Parameters.scala 47:9]
  wire  requestROI_4_0; // @[Parameters.scala 47:9]
  wire  requestROI_5_0; // @[Parameters.scala 47:9]
  wire  requestROI_6_0; // @[Parameters.scala 47:9]
  wire  requestROI_7_0; // @[Parameters.scala 47:9]
  wire  requestROI_8_0; // @[Parameters.scala 47:9]
  wire  requestROI_9_0; // @[Parameters.scala 47:9]
  wire  requestROI_10_0; // @[Parameters.scala 47:9]
  wire  requestROI_11_0; // @[Parameters.scala 47:9]
  wire  requestROI_12_0; // @[Parameters.scala 47:9]
  wire  requestBOI_0_0; // @[Parameters.scala 47:9]
  wire  requestBOI_1_0; // @[Parameters.scala 47:9]
  wire  requestBOI_2_0; // @[Parameters.scala 47:9]
  wire  requestBOI_3_0; // @[Parameters.scala 47:9]
  wire  requestBOI_4_0; // @[Parameters.scala 47:9]
  wire  requestBOI_5_0; // @[Parameters.scala 47:9]
  wire  requestBOI_6_0; // @[Parameters.scala 47:9]
  wire  requestBOI_7_0; // @[Parameters.scala 47:9]
  wire  requestBOI_8_0; // @[Parameters.scala 47:9]
  wire  requestBOI_9_0; // @[Parameters.scala 47:9]
  wire  requestBOI_10_0; // @[Parameters.scala 47:9]
  wire  requestBOI_11_0; // @[Parameters.scala 47:9]
  wire  requestBOI_12_0; // @[Parameters.scala 47:9]
  wire [5:0] _T_134; // @[Xbar.scala 64:75]
  wire [6:0] _T_140; // @[Xbar.scala 64:75]
  wire [12:0] _T_141; // @[Xbar.scala 64:75]
  wire  requestWIO_0_0; // @[Xbar.scala 65:73]
  wire  requestWIO_0_1; // @[Xbar.scala 65:73]
  wire  requestWIO_0_2; // @[Xbar.scala 65:73]
  wire  requestWIO_0_3; // @[Xbar.scala 65:73]
  wire  requestWIO_0_4; // @[Xbar.scala 65:73]
  wire  requestWIO_0_5; // @[Xbar.scala 65:73]
  wire  requestWIO_0_6; // @[Xbar.scala 65:73]
  wire  requestWIO_0_7; // @[Xbar.scala 65:73]
  wire  requestWIO_0_8; // @[Xbar.scala 65:73]
  wire  requestWIO_0_9; // @[Xbar.scala 65:73]
  wire  requestWIO_0_10; // @[Xbar.scala 65:73]
  wire  requestWIO_0_11; // @[Xbar.scala 65:73]
  wire  requestWIO_0_12; // @[Xbar.scala 65:73]
  wire [5:0] _T_152; // @[Xbar.scala 93:45]
  wire [12:0] _T_159; // @[Xbar.scala 93:45]
  wire  _T_162; // @[OneHot.scala 32:14]
  wire [7:0] _GEN_62; // @[OneHot.scala 32:28]
  wire [7:0] _T_163; // @[OneHot.scala 32:28]
  wire  _T_166; // @[OneHot.scala 32:14]
  wire [3:0] _T_167; // @[OneHot.scala 32:28]
  wire  _T_170; // @[OneHot.scala 32:14]
  wire [1:0] _T_171; // @[OneHot.scala 32:28]
  wire [3:0] _T_175; // @[Cat.scala 29:58]
  wire  _T_190; // @[OneHot.scala 32:14]
  wire [7:0] _GEN_63; // @[OneHot.scala 32:28]
  wire [7:0] _T_191; // @[OneHot.scala 32:28]
  wire  _T_194; // @[OneHot.scala 32:14]
  wire [3:0] _T_195; // @[OneHot.scala 32:28]
  wire  _T_198; // @[OneHot.scala 32:14]
  wire [1:0] _T_199; // @[OneHot.scala 32:28]
  wire [3:0] _T_203; // @[Cat.scala 29:58]
  wire  _T_292; // @[Mux.scala 27:72]
  wire  _T_293; // @[Mux.scala 27:72]
  wire  _T_305; // @[Mux.scala 27:72]
  wire  _T_294; // @[Mux.scala 27:72]
  wire  _T_306; // @[Mux.scala 27:72]
  wire  _T_295; // @[Mux.scala 27:72]
  wire  _T_307; // @[Mux.scala 27:72]
  wire  _T_296; // @[Mux.scala 27:72]
  wire  _T_308; // @[Mux.scala 27:72]
  wire  _T_297; // @[Mux.scala 27:72]
  wire  _T_309; // @[Mux.scala 27:72]
  wire  _T_298; // @[Mux.scala 27:72]
  wire  _T_310; // @[Mux.scala 27:72]
  wire  _T_299; // @[Mux.scala 27:72]
  wire  _T_311; // @[Mux.scala 27:72]
  wire  _T_300; // @[Mux.scala 27:72]
  wire  _T_312; // @[Mux.scala 27:72]
  wire  _T_301; // @[Mux.scala 27:72]
  wire  _T_313; // @[Mux.scala 27:72]
  wire  _T_302; // @[Mux.scala 27:72]
  wire  _T_314; // @[Mux.scala 27:72]
  wire  _T_303; // @[Mux.scala 27:72]
  wire  _T_315; // @[Mux.scala 27:72]
  wire  _T_304; // @[Mux.scala 27:72]
  wire  in_0_ar_ready; // @[Mux.scala 27:72]
  reg [2:0] _T_209; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_0;
  wire  _T_228; // @[Xbar.scala 112:22]
  reg [3:0] _T_210; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_1;
  wire  _T_227; // @[Xbar.scala 111:75]
  wire  _T_229; // @[Xbar.scala 112:34]
  wire  _T_230; // @[Xbar.scala 112:80]
  wire  _T_232; // @[Xbar.scala 112:48]
  wire  io_in_0_ar_ready; // @[Xbar.scala 130:45]
  wire  _T_204; // @[Decoupled.scala 40:37]
  reg  _T_1022; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_2;
  wire  _T_399; // @[Xbar.scala 222:40]
  wire  _T_401; // @[Xbar.scala 222:40]
  wire  _T_1023; // @[Xbar.scala 246:36]
  wire  _T_403; // @[Xbar.scala 222:40]
  wire  _T_1024; // @[Xbar.scala 246:36]
  wire  _T_405; // @[Xbar.scala 222:40]
  wire  _T_1025; // @[Xbar.scala 246:36]
  wire  _T_407; // @[Xbar.scala 222:40]
  wire  _T_1026; // @[Xbar.scala 246:36]
  wire  _T_409; // @[Xbar.scala 222:40]
  wire  _T_1027; // @[Xbar.scala 246:36]
  wire  _T_411; // @[Xbar.scala 222:40]
  wire  _T_1028; // @[Xbar.scala 246:36]
  wire  _T_413; // @[Xbar.scala 222:40]
  wire  _T_1029; // @[Xbar.scala 246:36]
  wire  _T_415; // @[Xbar.scala 222:40]
  wire  _T_1030; // @[Xbar.scala 246:36]
  wire  _T_417; // @[Xbar.scala 222:40]
  wire  _T_1031; // @[Xbar.scala 246:36]
  wire  _T_419; // @[Xbar.scala 222:40]
  wire  _T_1032; // @[Xbar.scala 246:36]
  wire  _T_421; // @[Xbar.scala 222:40]
  wire  _T_1033; // @[Xbar.scala 246:36]
  wire  _T_423; // @[Xbar.scala 222:40]
  wire  _T_1034; // @[Xbar.scala 246:36]
  reg  _T_1203_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_3;
  wire  _T_1220; // @[Mux.scala 27:72]
  reg  _T_1203_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_4;
  wire  _T_1221; // @[Mux.scala 27:72]
  wire  _T_1233; // @[Mux.scala 27:72]
  reg  _T_1203_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_5;
  wire  _T_1222; // @[Mux.scala 27:72]
  wire  _T_1234; // @[Mux.scala 27:72]
  reg  _T_1203_3; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_6;
  wire  _T_1223; // @[Mux.scala 27:72]
  wire  _T_1235; // @[Mux.scala 27:72]
  reg  _T_1203_4; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_7;
  wire  _T_1224; // @[Mux.scala 27:72]
  wire  _T_1236; // @[Mux.scala 27:72]
  reg  _T_1203_5; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_8;
  wire  _T_1225; // @[Mux.scala 27:72]
  wire  _T_1237; // @[Mux.scala 27:72]
  reg  _T_1203_6; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_9;
  wire  _T_1226; // @[Mux.scala 27:72]
  wire  _T_1238; // @[Mux.scala 27:72]
  reg  _T_1203_7; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_10;
  wire  _T_1227; // @[Mux.scala 27:72]
  wire  _T_1239; // @[Mux.scala 27:72]
  reg  _T_1203_8; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_11;
  wire  _T_1228; // @[Mux.scala 27:72]
  wire  _T_1240; // @[Mux.scala 27:72]
  reg  _T_1203_9; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_12;
  wire  _T_1229; // @[Mux.scala 27:72]
  wire  _T_1241; // @[Mux.scala 27:72]
  reg  _T_1203_10; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_13;
  wire  _T_1230; // @[Mux.scala 27:72]
  wire  _T_1242; // @[Mux.scala 27:72]
  reg  _T_1203_11; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_14;
  wire  _T_1231; // @[Mux.scala 27:72]
  wire  _T_1243; // @[Mux.scala 27:72]
  reg  _T_1203_12; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_15;
  wire  _T_1232; // @[Mux.scala 27:72]
  wire  _T_1244; // @[Mux.scala 27:72]
  wire  in_0_r_valid; // @[Xbar.scala 278:22]
  wire  _T_206; // @[Decoupled.scala 40:37]
  wire [5:0] _T_1039; // @[Cat.scala 29:58]
  wire [12:0] _T_1046; // @[Cat.scala 29:58]
  reg [12:0] _T_1053; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_16;
  wire [12:0] _T_1054; // @[Arbiter.scala 21:30]
  wire [12:0] _T_1055; // @[Arbiter.scala 21:28]
  wire [25:0] _T_1056; // @[Cat.scala 29:58]
  wire [25:0] _GEN_64; // @[package.scala 208:43]
  wire [25:0] _T_1058; // @[package.scala 208:43]
  wire [25:0] _GEN_65; // @[package.scala 208:43]
  wire [25:0] _T_1060; // @[package.scala 208:43]
  wire [25:0] _GEN_66; // @[package.scala 208:43]
  wire [25:0] _T_1062; // @[package.scala 208:43]
  wire [25:0] _GEN_67; // @[package.scala 208:43]
  wire [25:0] _T_1064; // @[package.scala 208:43]
  wire [25:0] _T_1067; // @[Arbiter.scala 22:66]
  wire [25:0] _GEN_68; // @[Arbiter.scala 22:58]
  wire [25:0] _T_1068; // @[Arbiter.scala 22:58]
  wire [12:0] _T_1071; // @[Arbiter.scala 23:39]
  wire [12:0] _T_1072; // @[Arbiter.scala 23:18]
  wire  _T_1104; // @[Xbar.scala 250:63]
  wire  _T_1204_0; // @[Xbar.scala 262:23]
  wire [35:0] _T_1249; // @[Mux.scala 27:72]
  wire [35:0] _T_1250; // @[Mux.scala 27:72]
  wire  _T_1105; // @[Xbar.scala 250:63]
  wire  _T_1204_1; // @[Xbar.scala 262:23]
  wire [35:0] _T_1253; // @[Mux.scala 27:72]
  wire [35:0] _T_1254; // @[Mux.scala 27:72]
  wire [35:0] _T_1299; // @[Mux.scala 27:72]
  wire  _T_1106; // @[Xbar.scala 250:63]
  wire  _T_1204_2; // @[Xbar.scala 262:23]
  wire [35:0] _T_1257; // @[Mux.scala 27:72]
  wire [35:0] _T_1258; // @[Mux.scala 27:72]
  wire [35:0] _T_1300; // @[Mux.scala 27:72]
  wire  _T_1107; // @[Xbar.scala 250:63]
  wire  _T_1204_3; // @[Xbar.scala 262:23]
  wire [35:0] _T_1261; // @[Mux.scala 27:72]
  wire [35:0] _T_1262; // @[Mux.scala 27:72]
  wire [35:0] _T_1301; // @[Mux.scala 27:72]
  wire  _T_1108; // @[Xbar.scala 250:63]
  wire  _T_1204_4; // @[Xbar.scala 262:23]
  wire [35:0] _T_1265; // @[Mux.scala 27:72]
  wire [35:0] _T_1266; // @[Mux.scala 27:72]
  wire [35:0] _T_1302; // @[Mux.scala 27:72]
  wire  _T_1109; // @[Xbar.scala 250:63]
  wire  _T_1204_5; // @[Xbar.scala 262:23]
  wire [35:0] _T_1269; // @[Mux.scala 27:72]
  wire [35:0] _T_1270; // @[Mux.scala 27:72]
  wire [35:0] _T_1303; // @[Mux.scala 27:72]
  wire  _T_1110; // @[Xbar.scala 250:63]
  wire  _T_1204_6; // @[Xbar.scala 262:23]
  wire [35:0] _T_1273; // @[Mux.scala 27:72]
  wire [35:0] _T_1274; // @[Mux.scala 27:72]
  wire [35:0] _T_1304; // @[Mux.scala 27:72]
  wire  _T_1111; // @[Xbar.scala 250:63]
  wire  _T_1204_7; // @[Xbar.scala 262:23]
  wire [35:0] _T_1277; // @[Mux.scala 27:72]
  wire [35:0] _T_1278; // @[Mux.scala 27:72]
  wire [35:0] _T_1305; // @[Mux.scala 27:72]
  wire  _T_1112; // @[Xbar.scala 250:63]
  wire  _T_1204_8; // @[Xbar.scala 262:23]
  wire [35:0] _T_1281; // @[Mux.scala 27:72]
  wire [35:0] _T_1282; // @[Mux.scala 27:72]
  wire [35:0] _T_1306; // @[Mux.scala 27:72]
  wire  _T_1113; // @[Xbar.scala 250:63]
  wire  _T_1204_9; // @[Xbar.scala 262:23]
  wire [35:0] _T_1285; // @[Mux.scala 27:72]
  wire [35:0] _T_1286; // @[Mux.scala 27:72]
  wire [35:0] _T_1307; // @[Mux.scala 27:72]
  wire  _T_1114; // @[Xbar.scala 250:63]
  wire  _T_1204_10; // @[Xbar.scala 262:23]
  wire [35:0] _T_1289; // @[Mux.scala 27:72]
  wire [35:0] _T_1290; // @[Mux.scala 27:72]
  wire [35:0] _T_1308; // @[Mux.scala 27:72]
  wire  _T_1115; // @[Xbar.scala 250:63]
  wire  _T_1204_11; // @[Xbar.scala 262:23]
  wire [35:0] _T_1293; // @[Mux.scala 27:72]
  wire [35:0] _T_1294; // @[Mux.scala 27:72]
  wire [35:0] _T_1309; // @[Mux.scala 27:72]
  wire  _T_1116; // @[Xbar.scala 250:63]
  wire  _T_1204_12; // @[Xbar.scala 262:23]
  wire [35:0] _T_1297; // @[Mux.scala 27:72]
  wire [35:0] _T_1298; // @[Mux.scala 27:72]
  wire [35:0] _T_1310; // @[Mux.scala 27:72]
  wire  in_0_r_bits_last; // @[Mux.scala 27:72]
  wire  _T_208; // @[Xbar.scala 120:45]
  wire [2:0] _GEN_69; // @[Xbar.scala 106:30]
  wire [2:0] _T_212; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_70; // @[Xbar.scala 106:48]
  wire [2:0] _T_214; // @[Xbar.scala 106:48]
  wire  _T_215; // @[Xbar.scala 107:23]
  wire  _T_216; // @[Xbar.scala 107:43]
  wire  _T_217; // @[Xbar.scala 107:34]
  wire  _T_219; // @[Xbar.scala 107:22]
  wire  _T_220; // @[Xbar.scala 107:22]
  wire  _T_221; // @[Xbar.scala 108:23]
  wire  _T_223; // @[Xbar.scala 108:34]
  wire  _T_225; // @[Xbar.scala 108:22]
  wire  _T_226; // @[Xbar.scala 108:22]
  wire  _T_332; // @[Mux.scala 27:72]
  wire  _T_333; // @[Mux.scala 27:72]
  wire  _T_345; // @[Mux.scala 27:72]
  wire  _T_334; // @[Mux.scala 27:72]
  wire  _T_346; // @[Mux.scala 27:72]
  wire  _T_335; // @[Mux.scala 27:72]
  wire  _T_347; // @[Mux.scala 27:72]
  wire  _T_336; // @[Mux.scala 27:72]
  wire  _T_348; // @[Mux.scala 27:72]
  wire  _T_337; // @[Mux.scala 27:72]
  wire  _T_349; // @[Mux.scala 27:72]
  wire  _T_338; // @[Mux.scala 27:72]
  wire  _T_350; // @[Mux.scala 27:72]
  wire  _T_339; // @[Mux.scala 27:72]
  wire  _T_351; // @[Mux.scala 27:72]
  wire  _T_340; // @[Mux.scala 27:72]
  wire  _T_352; // @[Mux.scala 27:72]
  wire  _T_341; // @[Mux.scala 27:72]
  wire  _T_353; // @[Mux.scala 27:72]
  wire  _T_342; // @[Mux.scala 27:72]
  wire  _T_354; // @[Mux.scala 27:72]
  wire  _T_343; // @[Mux.scala 27:72]
  wire  _T_355; // @[Mux.scala 27:72]
  wire  _T_344; // @[Mux.scala 27:72]
  wire  in_0_aw_ready; // @[Mux.scala 27:72]
  reg  _T_263; // @[Xbar.scala 137:30]
  reg [31:0] _RAND_17;
  wire  _T_267; // @[Xbar.scala 139:57]
  wire  _T_268; // @[Xbar.scala 139:45]
  reg [2:0] _T_237; // @[Xbar.scala 104:34]
  reg [31:0] _RAND_18;
  wire  _T_256; // @[Xbar.scala 112:22]
  reg [3:0] _T_238; // @[Xbar.scala 105:29]
  reg [31:0] _RAND_19;
  wire  _T_255; // @[Xbar.scala 111:75]
  wire  _T_257; // @[Xbar.scala 112:34]
  wire  _T_258; // @[Xbar.scala 112:80]
  wire  _T_260; // @[Xbar.scala 112:48]
  wire  io_in_0_aw_ready; // @[Xbar.scala 139:82]
  wire  _T_233; // @[Decoupled.scala 40:37]
  reg  _T_1317; // @[Xbar.scala 242:23]
  reg [31:0] _RAND_20;
  wire  _T_425; // @[Xbar.scala 222:40]
  wire  _T_427; // @[Xbar.scala 222:40]
  wire  _T_1318; // @[Xbar.scala 246:36]
  wire  _T_429; // @[Xbar.scala 222:40]
  wire  _T_1319; // @[Xbar.scala 246:36]
  wire  _T_431; // @[Xbar.scala 222:40]
  wire  _T_1320; // @[Xbar.scala 246:36]
  wire  _T_433; // @[Xbar.scala 222:40]
  wire  _T_1321; // @[Xbar.scala 246:36]
  wire  _T_435; // @[Xbar.scala 222:40]
  wire  _T_1322; // @[Xbar.scala 246:36]
  wire  _T_437; // @[Xbar.scala 222:40]
  wire  _T_1323; // @[Xbar.scala 246:36]
  wire  _T_439; // @[Xbar.scala 222:40]
  wire  _T_1324; // @[Xbar.scala 246:36]
  wire  _T_441; // @[Xbar.scala 222:40]
  wire  _T_1325; // @[Xbar.scala 246:36]
  wire  _T_443; // @[Xbar.scala 222:40]
  wire  _T_1326; // @[Xbar.scala 246:36]
  wire  _T_445; // @[Xbar.scala 222:40]
  wire  _T_1327; // @[Xbar.scala 246:36]
  wire  _T_447; // @[Xbar.scala 222:40]
  wire  _T_1328; // @[Xbar.scala 246:36]
  wire  _T_449; // @[Xbar.scala 222:40]
  wire  _T_1329; // @[Xbar.scala 246:36]
  reg  _T_1498_0; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_21;
  wire  _T_1515; // @[Mux.scala 27:72]
  reg  _T_1498_1; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_22;
  wire  _T_1516; // @[Mux.scala 27:72]
  wire  _T_1528; // @[Mux.scala 27:72]
  reg  _T_1498_2; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_23;
  wire  _T_1517; // @[Mux.scala 27:72]
  wire  _T_1529; // @[Mux.scala 27:72]
  reg  _T_1498_3; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_24;
  wire  _T_1518; // @[Mux.scala 27:72]
  wire  _T_1530; // @[Mux.scala 27:72]
  reg  _T_1498_4; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_25;
  wire  _T_1519; // @[Mux.scala 27:72]
  wire  _T_1531; // @[Mux.scala 27:72]
  reg  _T_1498_5; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_26;
  wire  _T_1520; // @[Mux.scala 27:72]
  wire  _T_1532; // @[Mux.scala 27:72]
  reg  _T_1498_6; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_27;
  wire  _T_1521; // @[Mux.scala 27:72]
  wire  _T_1533; // @[Mux.scala 27:72]
  reg  _T_1498_7; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_28;
  wire  _T_1522; // @[Mux.scala 27:72]
  wire  _T_1534; // @[Mux.scala 27:72]
  reg  _T_1498_8; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_29;
  wire  _T_1523; // @[Mux.scala 27:72]
  wire  _T_1535; // @[Mux.scala 27:72]
  reg  _T_1498_9; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_30;
  wire  _T_1524; // @[Mux.scala 27:72]
  wire  _T_1536; // @[Mux.scala 27:72]
  reg  _T_1498_10; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_31;
  wire  _T_1525; // @[Mux.scala 27:72]
  wire  _T_1537; // @[Mux.scala 27:72]
  reg  _T_1498_11; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_32;
  wire  _T_1526; // @[Mux.scala 27:72]
  wire  _T_1538; // @[Mux.scala 27:72]
  reg  _T_1498_12; // @[Xbar.scala 261:24]
  reg [31:0] _RAND_33;
  wire  _T_1527; // @[Mux.scala 27:72]
  wire  _T_1539; // @[Mux.scala 27:72]
  wire  in_0_b_valid; // @[Xbar.scala 278:22]
  wire  _T_235; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_71; // @[Xbar.scala 106:30]
  wire [2:0] _T_240; // @[Xbar.scala 106:30]
  wire [2:0] _GEN_72; // @[Xbar.scala 106:48]
  wire [2:0] _T_242; // @[Xbar.scala 106:48]
  wire  _T_243; // @[Xbar.scala 107:23]
  wire  _T_244; // @[Xbar.scala 107:43]
  wire  _T_245; // @[Xbar.scala 107:34]
  wire  _T_247; // @[Xbar.scala 107:22]
  wire  _T_248; // @[Xbar.scala 107:22]
  wire  _T_249; // @[Xbar.scala 108:23]
  wire  _T_251; // @[Xbar.scala 108:34]
  wire  _T_253; // @[Xbar.scala 108:22]
  wire  _T_254; // @[Xbar.scala 108:22]
  wire  in_0_ar_valid; // @[Xbar.scala 129:45]
  wire  _T_265; // @[Xbar.scala 138:45]
  wire  in_0_aw_valid; // @[Xbar.scala 138:82]
  wire  _T_270; // @[Xbar.scala 140:54]
  wire  _T_272; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[Xbar.scala 141:38]
  wire  _T_273; // @[Decoupled.scala 40:37]
  wire  in_0_w_valid; // @[Xbar.scala 145:43]
  wire  _T_372; // @[Mux.scala 27:72]
  wire  _T_373; // @[Mux.scala 27:72]
  wire  _T_385; // @[Mux.scala 27:72]
  wire  _T_374; // @[Mux.scala 27:72]
  wire  _T_386; // @[Mux.scala 27:72]
  wire  _T_375; // @[Mux.scala 27:72]
  wire  _T_387; // @[Mux.scala 27:72]
  wire  _T_376; // @[Mux.scala 27:72]
  wire  _T_388; // @[Mux.scala 27:72]
  wire  _T_377; // @[Mux.scala 27:72]
  wire  _T_389; // @[Mux.scala 27:72]
  wire  _T_378; // @[Mux.scala 27:72]
  wire  _T_390; // @[Mux.scala 27:72]
  wire  _T_379; // @[Mux.scala 27:72]
  wire  _T_391; // @[Mux.scala 27:72]
  wire  _T_380; // @[Mux.scala 27:72]
  wire  _T_392; // @[Mux.scala 27:72]
  wire  _T_381; // @[Mux.scala 27:72]
  wire  _T_393; // @[Mux.scala 27:72]
  wire  _T_382; // @[Mux.scala 27:72]
  wire  _T_394; // @[Mux.scala 27:72]
  wire  _T_383; // @[Mux.scala 27:72]
  wire  _T_395; // @[Mux.scala 27:72]
  wire  _T_384; // @[Mux.scala 27:72]
  wire  in_0_w_ready; // @[Mux.scala 27:72]
  wire  _T_276; // @[Xbar.scala 147:50]
  wire  out_0_ar_valid; // @[Xbar.scala 222:40]
  wire  out_1_ar_valid; // @[Xbar.scala 222:40]
  wire  out_2_ar_valid; // @[Xbar.scala 222:40]
  wire  out_3_ar_valid; // @[Xbar.scala 222:40]
  wire  out_4_ar_valid; // @[Xbar.scala 222:40]
  wire  out_5_ar_valid; // @[Xbar.scala 222:40]
  wire  out_6_ar_valid; // @[Xbar.scala 222:40]
  wire  out_7_ar_valid; // @[Xbar.scala 222:40]
  wire  out_8_ar_valid; // @[Xbar.scala 222:40]
  wire  out_9_ar_valid; // @[Xbar.scala 222:40]
  wire  out_10_ar_valid; // @[Xbar.scala 222:40]
  wire  out_11_ar_valid; // @[Xbar.scala 222:40]
  wire  out_12_ar_valid; // @[Xbar.scala 222:40]
  wire  out_0_aw_valid; // @[Xbar.scala 222:40]
  wire  out_1_aw_valid; // @[Xbar.scala 222:40]
  wire  out_2_aw_valid; // @[Xbar.scala 222:40]
  wire  out_3_aw_valid; // @[Xbar.scala 222:40]
  wire  out_4_aw_valid; // @[Xbar.scala 222:40]
  wire  out_5_aw_valid; // @[Xbar.scala 222:40]
  wire  out_6_aw_valid; // @[Xbar.scala 222:40]
  wire  out_7_aw_valid; // @[Xbar.scala 222:40]
  wire  out_8_aw_valid; // @[Xbar.scala 222:40]
  wire  out_9_aw_valid; // @[Xbar.scala 222:40]
  wire  out_10_aw_valid; // @[Xbar.scala 222:40]
  wire  out_11_aw_valid; // @[Xbar.scala 222:40]
  wire  out_12_aw_valid; // @[Xbar.scala 222:40]
  wire  _T_456; // @[Xbar.scala 256:60]
  wire  _T_462; // @[Xbar.scala 258:23]
  wire  _T_464; // @[Xbar.scala 258:12]
  wire  _T_465; // @[Xbar.scala 258:12]
  wire  _T_477; // @[Xbar.scala 256:60]
  wire  _T_483; // @[Xbar.scala 258:23]
  wire  _T_485; // @[Xbar.scala 258:12]
  wire  _T_486; // @[Xbar.scala 258:12]
  wire  _T_500; // @[Xbar.scala 256:60]
  wire  _T_506; // @[Xbar.scala 258:23]
  wire  _T_508; // @[Xbar.scala 258:12]
  wire  _T_509; // @[Xbar.scala 258:12]
  wire  _T_521; // @[Xbar.scala 256:60]
  wire  _T_527; // @[Xbar.scala 258:23]
  wire  _T_529; // @[Xbar.scala 258:12]
  wire  _T_530; // @[Xbar.scala 258:12]
  wire  _T_544; // @[Xbar.scala 256:60]
  wire  _T_550; // @[Xbar.scala 258:23]
  wire  _T_552; // @[Xbar.scala 258:12]
  wire  _T_553; // @[Xbar.scala 258:12]
  wire  _T_565; // @[Xbar.scala 256:60]
  wire  _T_571; // @[Xbar.scala 258:23]
  wire  _T_573; // @[Xbar.scala 258:12]
  wire  _T_574; // @[Xbar.scala 258:12]
  wire  _T_588; // @[Xbar.scala 256:60]
  wire  _T_594; // @[Xbar.scala 258:23]
  wire  _T_596; // @[Xbar.scala 258:12]
  wire  _T_597; // @[Xbar.scala 258:12]
  wire  _T_609; // @[Xbar.scala 256:60]
  wire  _T_615; // @[Xbar.scala 258:23]
  wire  _T_617; // @[Xbar.scala 258:12]
  wire  _T_618; // @[Xbar.scala 258:12]
  wire  _T_632; // @[Xbar.scala 256:60]
  wire  _T_638; // @[Xbar.scala 258:23]
  wire  _T_640; // @[Xbar.scala 258:12]
  wire  _T_641; // @[Xbar.scala 258:12]
  wire  _T_653; // @[Xbar.scala 256:60]
  wire  _T_659; // @[Xbar.scala 258:23]
  wire  _T_661; // @[Xbar.scala 258:12]
  wire  _T_662; // @[Xbar.scala 258:12]
  wire  _T_676; // @[Xbar.scala 256:60]
  wire  _T_682; // @[Xbar.scala 258:23]
  wire  _T_684; // @[Xbar.scala 258:12]
  wire  _T_685; // @[Xbar.scala 258:12]
  wire  _T_697; // @[Xbar.scala 256:60]
  wire  _T_703; // @[Xbar.scala 258:23]
  wire  _T_705; // @[Xbar.scala 258:12]
  wire  _T_706; // @[Xbar.scala 258:12]
  wire  _T_720; // @[Xbar.scala 256:60]
  wire  _T_726; // @[Xbar.scala 258:23]
  wire  _T_728; // @[Xbar.scala 258:12]
  wire  _T_729; // @[Xbar.scala 258:12]
  wire  _T_741; // @[Xbar.scala 256:60]
  wire  _T_747; // @[Xbar.scala 258:23]
  wire  _T_749; // @[Xbar.scala 258:12]
  wire  _T_750; // @[Xbar.scala 258:12]
  wire  _T_764; // @[Xbar.scala 256:60]
  wire  _T_770; // @[Xbar.scala 258:23]
  wire  _T_772; // @[Xbar.scala 258:12]
  wire  _T_773; // @[Xbar.scala 258:12]
  wire  _T_785; // @[Xbar.scala 256:60]
  wire  _T_791; // @[Xbar.scala 258:23]
  wire  _T_793; // @[Xbar.scala 258:12]
  wire  _T_794; // @[Xbar.scala 258:12]
  wire  _T_808; // @[Xbar.scala 256:60]
  wire  _T_814; // @[Xbar.scala 258:23]
  wire  _T_816; // @[Xbar.scala 258:12]
  wire  _T_817; // @[Xbar.scala 258:12]
  wire  _T_829; // @[Xbar.scala 256:60]
  wire  _T_835; // @[Xbar.scala 258:23]
  wire  _T_837; // @[Xbar.scala 258:12]
  wire  _T_838; // @[Xbar.scala 258:12]
  wire  _T_852; // @[Xbar.scala 256:60]
  wire  _T_858; // @[Xbar.scala 258:23]
  wire  _T_860; // @[Xbar.scala 258:12]
  wire  _T_861; // @[Xbar.scala 258:12]
  wire  _T_873; // @[Xbar.scala 256:60]
  wire  _T_879; // @[Xbar.scala 258:23]
  wire  _T_881; // @[Xbar.scala 258:12]
  wire  _T_882; // @[Xbar.scala 258:12]
  wire  _T_896; // @[Xbar.scala 256:60]
  wire  _T_902; // @[Xbar.scala 258:23]
  wire  _T_904; // @[Xbar.scala 258:12]
  wire  _T_905; // @[Xbar.scala 258:12]
  wire  _T_917; // @[Xbar.scala 256:60]
  wire  _T_923; // @[Xbar.scala 258:23]
  wire  _T_925; // @[Xbar.scala 258:12]
  wire  _T_926; // @[Xbar.scala 258:12]
  wire  _T_940; // @[Xbar.scala 256:60]
  wire  _T_946; // @[Xbar.scala 258:23]
  wire  _T_948; // @[Xbar.scala 258:12]
  wire  _T_949; // @[Xbar.scala 258:12]
  wire  _T_961; // @[Xbar.scala 256:60]
  wire  _T_967; // @[Xbar.scala 258:23]
  wire  _T_969; // @[Xbar.scala 258:12]
  wire  _T_970; // @[Xbar.scala 258:12]
  wire  _T_984; // @[Xbar.scala 256:60]
  wire  _T_990; // @[Xbar.scala 258:23]
  wire  _T_992; // @[Xbar.scala 258:12]
  wire  _T_993; // @[Xbar.scala 258:12]
  wire  _T_1005; // @[Xbar.scala 256:60]
  wire  _T_1011; // @[Xbar.scala 258:23]
  wire  _T_1013; // @[Xbar.scala 258:12]
  wire  _T_1014; // @[Xbar.scala 258:12]
  wire  _T_1073; // @[Arbiter.scala 24:27]
  wire  _T_1074; // @[Arbiter.scala 24:18]
  wire [12:0] _T_1075; // @[Arbiter.scala 25:29]
  wire [13:0] _T_1076; // @[package.scala 199:48]
  wire [12:0] _T_1078; // @[package.scala 199:43]
  wire [14:0] _T_1079; // @[package.scala 199:48]
  wire [12:0] _T_1081; // @[package.scala 199:43]
  wire [16:0] _T_1082; // @[package.scala 199:48]
  wire [12:0] _T_1084; // @[package.scala 199:43]
  wire [20:0] _T_1085; // @[package.scala 199:48]
  wire [12:0] _T_1087; // @[package.scala 199:43]
  wire  _T_1119; // @[Xbar.scala 255:50]
  wire  _T_1120; // @[Xbar.scala 255:50]
  wire  _T_1121; // @[Xbar.scala 255:50]
  wire  _T_1122; // @[Xbar.scala 255:50]
  wire  _T_1123; // @[Xbar.scala 255:50]
  wire  _T_1124; // @[Xbar.scala 255:50]
  wire  _T_1125; // @[Xbar.scala 255:50]
  wire  _T_1126; // @[Xbar.scala 255:50]
  wire  _T_1127; // @[Xbar.scala 255:50]
  wire  _T_1128; // @[Xbar.scala 255:50]
  wire  _T_1129; // @[Xbar.scala 255:50]
  wire  _T_1130; // @[Xbar.scala 255:50]
  wire  _T_1132; // @[Xbar.scala 256:60]
  wire  _T_1135; // @[Xbar.scala 256:60]
  wire  _T_1136; // @[Xbar.scala 256:57]
  wire  _T_1137; // @[Xbar.scala 256:54]
  wire  _T_1138; // @[Xbar.scala 256:60]
  wire  _T_1139; // @[Xbar.scala 256:57]
  wire  _T_1140; // @[Xbar.scala 256:54]
  wire  _T_1141; // @[Xbar.scala 256:60]
  wire  _T_1142; // @[Xbar.scala 256:57]
  wire  _T_1143; // @[Xbar.scala 256:54]
  wire  _T_1144; // @[Xbar.scala 256:60]
  wire  _T_1145; // @[Xbar.scala 256:57]
  wire  _T_1146; // @[Xbar.scala 256:54]
  wire  _T_1147; // @[Xbar.scala 256:60]
  wire  _T_1148; // @[Xbar.scala 256:57]
  wire  _T_1149; // @[Xbar.scala 256:54]
  wire  _T_1150; // @[Xbar.scala 256:60]
  wire  _T_1151; // @[Xbar.scala 256:57]
  wire  _T_1152; // @[Xbar.scala 256:54]
  wire  _T_1153; // @[Xbar.scala 256:60]
  wire  _T_1154; // @[Xbar.scala 256:57]
  wire  _T_1155; // @[Xbar.scala 256:54]
  wire  _T_1156; // @[Xbar.scala 256:60]
  wire  _T_1157; // @[Xbar.scala 256:57]
  wire  _T_1158; // @[Xbar.scala 256:54]
  wire  _T_1159; // @[Xbar.scala 256:60]
  wire  _T_1160; // @[Xbar.scala 256:57]
  wire  _T_1161; // @[Xbar.scala 256:54]
  wire  _T_1162; // @[Xbar.scala 256:60]
  wire  _T_1163; // @[Xbar.scala 256:57]
  wire  _T_1164; // @[Xbar.scala 256:54]
  wire  _T_1165; // @[Xbar.scala 256:60]
  wire  _T_1166; // @[Xbar.scala 256:57]
  wire  _T_1167; // @[Xbar.scala 256:54]
  wire  _T_1168; // @[Xbar.scala 256:60]
  wire  _T_1169; // @[Xbar.scala 256:57]
  wire  _T_1171; // @[Xbar.scala 256:75]
  wire  _T_1172; // @[Xbar.scala 256:75]
  wire  _T_1173; // @[Xbar.scala 256:75]
  wire  _T_1174; // @[Xbar.scala 256:75]
  wire  _T_1175; // @[Xbar.scala 256:75]
  wire  _T_1176; // @[Xbar.scala 256:75]
  wire  _T_1177; // @[Xbar.scala 256:75]
  wire  _T_1178; // @[Xbar.scala 256:75]
  wire  _T_1179; // @[Xbar.scala 256:75]
  wire  _T_1180; // @[Xbar.scala 256:75]
  wire  _T_1181; // @[Xbar.scala 256:75]
  wire  _T_1183; // @[Xbar.scala 256:11]
  wire  _T_1184; // @[Xbar.scala 256:11]
  wire  _T_1185; // @[Xbar.scala 258:13]
  wire  _T_1198; // @[Xbar.scala 258:23]
  wire  _T_1200; // @[Xbar.scala 258:12]
  wire  _T_1201; // @[Xbar.scala 258:12]
  wire  _GEN_57; // @[Xbar.scala 266:21]
  wire  _GEN_58; // @[Xbar.scala 267:24]
  wire  _T_1206_0; // @[Xbar.scala 270:24]
  wire  _T_1206_1; // @[Xbar.scala 270:24]
  wire  _T_1206_2; // @[Xbar.scala 270:24]
  wire  _T_1206_3; // @[Xbar.scala 270:24]
  wire  _T_1206_4; // @[Xbar.scala 270:24]
  wire  _T_1206_5; // @[Xbar.scala 270:24]
  wire  _T_1206_6; // @[Xbar.scala 270:24]
  wire  _T_1206_7; // @[Xbar.scala 270:24]
  wire  _T_1206_8; // @[Xbar.scala 270:24]
  wire  _T_1206_9; // @[Xbar.scala 270:24]
  wire  _T_1206_10; // @[Xbar.scala 270:24]
  wire  _T_1206_11; // @[Xbar.scala 270:24]
  wire  _T_1206_12; // @[Xbar.scala 270:24]
  wire [5:0] _T_1334; // @[Cat.scala 29:58]
  wire [12:0] _T_1341; // @[Cat.scala 29:58]
  reg [12:0] _T_1348; // @[Arbiter.scala 20:23]
  reg [31:0] _RAND_34;
  wire [12:0] _T_1349; // @[Arbiter.scala 21:30]
  wire [12:0] _T_1350; // @[Arbiter.scala 21:28]
  wire [25:0] _T_1351; // @[Cat.scala 29:58]
  wire [25:0] _GEN_73; // @[package.scala 208:43]
  wire [25:0] _T_1353; // @[package.scala 208:43]
  wire [25:0] _GEN_74; // @[package.scala 208:43]
  wire [25:0] _T_1355; // @[package.scala 208:43]
  wire [25:0] _GEN_75; // @[package.scala 208:43]
  wire [25:0] _T_1357; // @[package.scala 208:43]
  wire [25:0] _GEN_76; // @[package.scala 208:43]
  wire [25:0] _T_1359; // @[package.scala 208:43]
  wire [25:0] _T_1362; // @[Arbiter.scala 22:66]
  wire [25:0] _GEN_77; // @[Arbiter.scala 22:58]
  wire [25:0] _T_1363; // @[Arbiter.scala 22:58]
  wire [12:0] _T_1366; // @[Arbiter.scala 23:39]
  wire [12:0] _T_1367; // @[Arbiter.scala 23:18]
  wire  _T_1368; // @[Arbiter.scala 24:27]
  wire  _T_1369; // @[Arbiter.scala 24:18]
  wire [12:0] _T_1370; // @[Arbiter.scala 25:29]
  wire [13:0] _T_1371; // @[package.scala 199:48]
  wire [12:0] _T_1373; // @[package.scala 199:43]
  wire [14:0] _T_1374; // @[package.scala 199:48]
  wire [12:0] _T_1376; // @[package.scala 199:43]
  wire [16:0] _T_1377; // @[package.scala 199:48]
  wire [12:0] _T_1379; // @[package.scala 199:43]
  wire [20:0] _T_1380; // @[package.scala 199:48]
  wire [12:0] _T_1382; // @[package.scala 199:43]
  wire  _T_1399; // @[Xbar.scala 250:63]
  wire  _T_1400; // @[Xbar.scala 250:63]
  wire  _T_1401; // @[Xbar.scala 250:63]
  wire  _T_1402; // @[Xbar.scala 250:63]
  wire  _T_1403; // @[Xbar.scala 250:63]
  wire  _T_1404; // @[Xbar.scala 250:63]
  wire  _T_1405; // @[Xbar.scala 250:63]
  wire  _T_1406; // @[Xbar.scala 250:63]
  wire  _T_1407; // @[Xbar.scala 250:63]
  wire  _T_1408; // @[Xbar.scala 250:63]
  wire  _T_1409; // @[Xbar.scala 250:63]
  wire  _T_1410; // @[Xbar.scala 250:63]
  wire  _T_1411; // @[Xbar.scala 250:63]
  wire  _T_1414; // @[Xbar.scala 255:50]
  wire  _T_1415; // @[Xbar.scala 255:50]
  wire  _T_1416; // @[Xbar.scala 255:50]
  wire  _T_1417; // @[Xbar.scala 255:50]
  wire  _T_1418; // @[Xbar.scala 255:50]
  wire  _T_1419; // @[Xbar.scala 255:50]
  wire  _T_1420; // @[Xbar.scala 255:50]
  wire  _T_1421; // @[Xbar.scala 255:50]
  wire  _T_1422; // @[Xbar.scala 255:50]
  wire  _T_1423; // @[Xbar.scala 255:50]
  wire  _T_1424; // @[Xbar.scala 255:50]
  wire  _T_1425; // @[Xbar.scala 255:50]
  wire  _T_1427; // @[Xbar.scala 256:60]
  wire  _T_1430; // @[Xbar.scala 256:60]
  wire  _T_1431; // @[Xbar.scala 256:57]
  wire  _T_1432; // @[Xbar.scala 256:54]
  wire  _T_1433; // @[Xbar.scala 256:60]
  wire  _T_1434; // @[Xbar.scala 256:57]
  wire  _T_1435; // @[Xbar.scala 256:54]
  wire  _T_1436; // @[Xbar.scala 256:60]
  wire  _T_1437; // @[Xbar.scala 256:57]
  wire  _T_1438; // @[Xbar.scala 256:54]
  wire  _T_1439; // @[Xbar.scala 256:60]
  wire  _T_1440; // @[Xbar.scala 256:57]
  wire  _T_1441; // @[Xbar.scala 256:54]
  wire  _T_1442; // @[Xbar.scala 256:60]
  wire  _T_1443; // @[Xbar.scala 256:57]
  wire  _T_1444; // @[Xbar.scala 256:54]
  wire  _T_1445; // @[Xbar.scala 256:60]
  wire  _T_1446; // @[Xbar.scala 256:57]
  wire  _T_1447; // @[Xbar.scala 256:54]
  wire  _T_1448; // @[Xbar.scala 256:60]
  wire  _T_1449; // @[Xbar.scala 256:57]
  wire  _T_1450; // @[Xbar.scala 256:54]
  wire  _T_1451; // @[Xbar.scala 256:60]
  wire  _T_1452; // @[Xbar.scala 256:57]
  wire  _T_1453; // @[Xbar.scala 256:54]
  wire  _T_1454; // @[Xbar.scala 256:60]
  wire  _T_1455; // @[Xbar.scala 256:57]
  wire  _T_1456; // @[Xbar.scala 256:54]
  wire  _T_1457; // @[Xbar.scala 256:60]
  wire  _T_1458; // @[Xbar.scala 256:57]
  wire  _T_1459; // @[Xbar.scala 256:54]
  wire  _T_1460; // @[Xbar.scala 256:60]
  wire  _T_1461; // @[Xbar.scala 256:57]
  wire  _T_1462; // @[Xbar.scala 256:54]
  wire  _T_1463; // @[Xbar.scala 256:60]
  wire  _T_1464; // @[Xbar.scala 256:57]
  wire  _T_1466; // @[Xbar.scala 256:75]
  wire  _T_1467; // @[Xbar.scala 256:75]
  wire  _T_1468; // @[Xbar.scala 256:75]
  wire  _T_1469; // @[Xbar.scala 256:75]
  wire  _T_1470; // @[Xbar.scala 256:75]
  wire  _T_1471; // @[Xbar.scala 256:75]
  wire  _T_1472; // @[Xbar.scala 256:75]
  wire  _T_1473; // @[Xbar.scala 256:75]
  wire  _T_1474; // @[Xbar.scala 256:75]
  wire  _T_1475; // @[Xbar.scala 256:75]
  wire  _T_1476; // @[Xbar.scala 256:75]
  wire  _T_1478; // @[Xbar.scala 256:11]
  wire  _T_1479; // @[Xbar.scala 256:11]
  wire  _T_1480; // @[Xbar.scala 258:13]
  wire  _T_1493; // @[Xbar.scala 258:23]
  wire  _T_1495; // @[Xbar.scala 258:12]
  wire  _T_1496; // @[Xbar.scala 258:12]
  wire  _T_1499_0; // @[Xbar.scala 262:23]
  wire  _T_1499_1; // @[Xbar.scala 262:23]
  wire  _T_1499_2; // @[Xbar.scala 262:23]
  wire  _T_1499_3; // @[Xbar.scala 262:23]
  wire  _T_1499_4; // @[Xbar.scala 262:23]
  wire  _T_1499_5; // @[Xbar.scala 262:23]
  wire  _T_1499_6; // @[Xbar.scala 262:23]
  wire  _T_1499_7; // @[Xbar.scala 262:23]
  wire  _T_1499_8; // @[Xbar.scala 262:23]
  wire  _T_1499_9; // @[Xbar.scala 262:23]
  wire  _T_1499_10; // @[Xbar.scala 262:23]
  wire  _T_1499_11; // @[Xbar.scala 262:23]
  wire  _T_1499_12; // @[Xbar.scala 262:23]
  wire  _GEN_60; // @[Xbar.scala 266:21]
  wire  _GEN_61; // @[Xbar.scala 267:24]
  wire  _T_1501_0; // @[Xbar.scala 270:24]
  wire  _T_1501_1; // @[Xbar.scala 270:24]
  wire  _T_1501_2; // @[Xbar.scala 270:24]
  wire  _T_1501_3; // @[Xbar.scala 270:24]
  wire  _T_1501_4; // @[Xbar.scala 270:24]
  wire  _T_1501_5; // @[Xbar.scala 270:24]
  wire  _T_1501_6; // @[Xbar.scala 270:24]
  wire  _T_1501_7; // @[Xbar.scala 270:24]
  wire  _T_1501_8; // @[Xbar.scala 270:24]
  wire  _T_1501_9; // @[Xbar.scala 270:24]
  wire  _T_1501_10; // @[Xbar.scala 270:24]
  wire  _T_1501_11; // @[Xbar.scala 270:24]
  wire  _T_1501_12; // @[Xbar.scala 270:24]
  wire [2:0] _T_1542; // @[Mux.scala 27:72]
  wire [2:0] _T_1543; // @[Mux.scala 27:72]
  wire [2:0] _T_1544; // @[Mux.scala 27:72]
  wire [2:0] _T_1545; // @[Mux.scala 27:72]
  wire [2:0] _T_1546; // @[Mux.scala 27:72]
  wire [2:0] _T_1547; // @[Mux.scala 27:72]
  wire [2:0] _T_1548; // @[Mux.scala 27:72]
  wire [2:0] _T_1549; // @[Mux.scala 27:72]
  wire [2:0] _T_1550; // @[Mux.scala 27:72]
  wire [2:0] _T_1551; // @[Mux.scala 27:72]
  wire [2:0] _T_1552; // @[Mux.scala 27:72]
  wire [2:0] _T_1553; // @[Mux.scala 27:72]
  wire [2:0] _T_1554; // @[Mux.scala 27:72]
  wire [2:0] _T_1555; // @[Mux.scala 27:72]
  wire [2:0] _T_1556; // @[Mux.scala 27:72]
  wire [2:0] _T_1557; // @[Mux.scala 27:72]
  wire [2:0] _T_1558; // @[Mux.scala 27:72]
  wire [2:0] _T_1559; // @[Mux.scala 27:72]
  wire [2:0] _T_1560; // @[Mux.scala 27:72]
  wire [2:0] _T_1561; // @[Mux.scala 27:72]
  wire [2:0] _T_1562; // @[Mux.scala 27:72]
  wire [2:0] _T_1563; // @[Mux.scala 27:72]
  wire [2:0] _T_1564; // @[Mux.scala 27:72]
  wire [2:0] _T_1565; // @[Mux.scala 27:72]
  wire [2:0] _T_1566; // @[Mux.scala 27:72]
  wire [2:0] _T_1567; // @[Mux.scala 27:72]
  wire [2:0] _T_1568; // @[Mux.scala 27:72]
  wire [2:0] _T_1569; // @[Mux.scala 27:72]
  wire [2:0] _T_1570; // @[Mux.scala 27:72]
  wire [2:0] _T_1571; // @[Mux.scala 27:72]
  wire [2:0] _T_1572; // @[Mux.scala 27:72]
  wire [2:0] _T_1573; // @[Mux.scala 27:72]
  wire [2:0] _T_1574; // @[Mux.scala 27:72]
  wire [2:0] _T_1575; // @[Mux.scala 27:72]
  wire [2:0] _T_1576; // @[Mux.scala 27:72]
  wire [2:0] _T_1577; // @[Mux.scala 27:72]
  wire [2:0] _T_1578; // @[Mux.scala 27:72]
  wire [2:0] _T_1579; // @[Mux.scala 27:72]
  QueueCompatibility_2 awIn_0 ( // @[Xbar.scala 55:47]
    .clock(awIn_0_clock),
    .reset(awIn_0_reset),
    .io_enq_ready(awIn_0_io_enq_ready),
    .io_enq_valid(awIn_0_io_enq_valid),
    .io_enq_bits(awIn_0_io_enq_bits),
    .io_deq_ready(awIn_0_io_deq_ready),
    .io_deq_valid(awIn_0_io_deq_valid),
    .io_deq_bits(awIn_0_io_deq_bits)
  );
  assign _T_1 = {1'b0,$signed(auto_in_ar_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_3 = $signed(_T_1) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_0 = $signed(_T_3) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_5 = auto_in_ar_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  assign _T_6 = {1'b0,$signed(_T_5)}; // @[Parameters.scala 137:49]
  assign _T_8 = $signed(_T_6) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestARIO_0_1 = $signed(_T_8) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_10 = auto_in_ar_bits_addr ^ 30'h1100; // @[Parameters.scala 137:31]
  assign _T_11 = {1'b0,$signed(_T_10)}; // @[Parameters.scala 137:49]
  assign _T_13 = $signed(_T_11) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_2 = $signed(_T_13) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_15 = auto_in_ar_bits_addr ^ 30'h3000; // @[Parameters.scala 137:31]
  assign _T_16 = {1'b0,$signed(_T_15)}; // @[Parameters.scala 137:49]
  assign _T_18 = $signed(_T_16) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestARIO_0_3 = $signed(_T_18) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_20 = auto_in_ar_bits_addr ^ 30'h3100; // @[Parameters.scala 137:31]
  assign _T_21 = {1'b0,$signed(_T_20)}; // @[Parameters.scala 137:49]
  assign _T_23 = $signed(_T_21) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_4 = $signed(_T_23) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_25 = auto_in_ar_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  assign _T_26 = {1'b0,$signed(_T_25)}; // @[Parameters.scala 137:49]
  assign _T_28 = $signed(_T_26) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestARIO_0_5 = $signed(_T_28) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_30 = auto_in_ar_bits_addr ^ 30'h2100; // @[Parameters.scala 137:31]
  assign _T_31 = {1'b0,$signed(_T_30)}; // @[Parameters.scala 137:49]
  assign _T_33 = $signed(_T_31) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_6 = $signed(_T_33) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_35 = auto_in_ar_bits_addr ^ 30'h4000; // @[Parameters.scala 137:31]
  assign _T_36 = {1'b0,$signed(_T_35)}; // @[Parameters.scala 137:49]
  assign _T_38 = $signed(_T_36) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestARIO_0_7 = $signed(_T_38) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_40 = auto_in_ar_bits_addr ^ 30'h4100; // @[Parameters.scala 137:31]
  assign _T_41 = {1'b0,$signed(_T_40)}; // @[Parameters.scala 137:49]
  assign _T_43 = $signed(_T_41) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_8 = $signed(_T_43) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_45 = auto_in_ar_bits_addr ^ 30'h5000; // @[Parameters.scala 137:31]
  assign _T_46 = {1'b0,$signed(_T_45)}; // @[Parameters.scala 137:49]
  assign _T_48 = $signed(_T_46) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_9 = $signed(_T_48) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_50 = auto_in_ar_bits_addr ^ 30'h5010; // @[Parameters.scala 137:31]
  assign _T_51 = {1'b0,$signed(_T_50)}; // @[Parameters.scala 137:49]
  assign _T_53 = $signed(_T_51) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_10 = $signed(_T_53) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_55 = auto_in_ar_bits_addr ^ 30'h6000; // @[Parameters.scala 137:31]
  assign _T_56 = {1'b0,$signed(_T_55)}; // @[Parameters.scala 137:49]
  assign _T_58 = $signed(_T_56) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestARIO_0_11 = $signed(_T_58) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_60 = auto_in_ar_bits_addr ^ 30'h6100; // @[Parameters.scala 137:31]
  assign _T_61 = {1'b0,$signed(_T_60)}; // @[Parameters.scala 137:49]
  assign _T_63 = $signed(_T_61) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestARIO_0_12 = $signed(_T_63) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_66 = {1'b0,$signed(auto_in_aw_bits_addr)}; // @[Parameters.scala 137:49]
  assign _T_68 = $signed(_T_66) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_0 = $signed(_T_68) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_70 = auto_in_aw_bits_addr ^ 30'h1000; // @[Parameters.scala 137:31]
  assign _T_71 = {1'b0,$signed(_T_70)}; // @[Parameters.scala 137:49]
  assign _T_73 = $signed(_T_71) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_1 = $signed(_T_73) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_75 = auto_in_aw_bits_addr ^ 30'h1100; // @[Parameters.scala 137:31]
  assign _T_76 = {1'b0,$signed(_T_75)}; // @[Parameters.scala 137:49]
  assign _T_78 = $signed(_T_76) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_2 = $signed(_T_78) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_80 = auto_in_aw_bits_addr ^ 30'h3000; // @[Parameters.scala 137:31]
  assign _T_81 = {1'b0,$signed(_T_80)}; // @[Parameters.scala 137:49]
  assign _T_83 = $signed(_T_81) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_3 = $signed(_T_83) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_85 = auto_in_aw_bits_addr ^ 30'h3100; // @[Parameters.scala 137:31]
  assign _T_86 = {1'b0,$signed(_T_85)}; // @[Parameters.scala 137:49]
  assign _T_88 = $signed(_T_86) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_4 = $signed(_T_88) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_90 = auto_in_aw_bits_addr ^ 30'h2000; // @[Parameters.scala 137:31]
  assign _T_91 = {1'b0,$signed(_T_90)}; // @[Parameters.scala 137:49]
  assign _T_93 = $signed(_T_91) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_5 = $signed(_T_93) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_95 = auto_in_aw_bits_addr ^ 30'h2100; // @[Parameters.scala 137:31]
  assign _T_96 = {1'b0,$signed(_T_95)}; // @[Parameters.scala 137:49]
  assign _T_98 = $signed(_T_96) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_6 = $signed(_T_98) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_100 = auto_in_aw_bits_addr ^ 30'h4000; // @[Parameters.scala 137:31]
  assign _T_101 = {1'b0,$signed(_T_100)}; // @[Parameters.scala 137:49]
  assign _T_103 = $signed(_T_101) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_7 = $signed(_T_103) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_105 = auto_in_aw_bits_addr ^ 30'h4100; // @[Parameters.scala 137:31]
  assign _T_106 = {1'b0,$signed(_T_105)}; // @[Parameters.scala 137:49]
  assign _T_108 = $signed(_T_106) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_8 = $signed(_T_108) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_110 = auto_in_aw_bits_addr ^ 30'h5000; // @[Parameters.scala 137:31]
  assign _T_111 = {1'b0,$signed(_T_110)}; // @[Parameters.scala 137:49]
  assign _T_113 = $signed(_T_111) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_9 = $signed(_T_113) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_115 = auto_in_aw_bits_addr ^ 30'h5010; // @[Parameters.scala 137:31]
  assign _T_116 = {1'b0,$signed(_T_115)}; // @[Parameters.scala 137:49]
  assign _T_118 = $signed(_T_116) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_10 = $signed(_T_118) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_120 = auto_in_aw_bits_addr ^ 30'h6000; // @[Parameters.scala 137:31]
  assign _T_121 = {1'b0,$signed(_T_120)}; // @[Parameters.scala 137:49]
  assign _T_123 = $signed(_T_121) & 31'sh7100; // @[Parameters.scala 137:52]
  assign requestAWIO_0_11 = $signed(_T_123) == 31'sh0; // @[Parameters.scala 137:67]
  assign _T_125 = auto_in_aw_bits_addr ^ 30'h6100; // @[Parameters.scala 137:31]
  assign _T_126 = {1'b0,$signed(_T_125)}; // @[Parameters.scala 137:49]
  assign _T_128 = $signed(_T_126) & 31'sh7110; // @[Parameters.scala 137:52]
  assign requestAWIO_0_12 = $signed(_T_128) == 31'sh0; // @[Parameters.scala 137:67]
  assign requestROI_0_0 = ~auto_out_0_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_1_0 = ~auto_out_1_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_2_0 = ~auto_out_2_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_3_0 = ~auto_out_3_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_4_0 = ~auto_out_4_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_5_0 = ~auto_out_5_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_6_0 = ~auto_out_6_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_7_0 = ~auto_out_7_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_8_0 = ~auto_out_8_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_9_0 = ~auto_out_9_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_10_0 = ~auto_out_10_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_11_0 = ~auto_out_11_r_bits_id; // @[Parameters.scala 47:9]
  assign requestROI_12_0 = ~auto_out_12_r_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_0_0 = ~auto_out_0_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_1_0 = ~auto_out_1_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_2_0 = ~auto_out_2_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_3_0 = ~auto_out_3_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_4_0 = ~auto_out_4_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_5_0 = ~auto_out_5_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_6_0 = ~auto_out_6_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_7_0 = ~auto_out_7_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_8_0 = ~auto_out_8_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_9_0 = ~auto_out_9_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_10_0 = ~auto_out_10_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_11_0 = ~auto_out_11_b_bits_id; // @[Parameters.scala 47:9]
  assign requestBOI_12_0 = ~auto_out_12_b_bits_id; // @[Parameters.scala 47:9]
  assign _T_134 = {requestAWIO_0_5,requestAWIO_0_4,requestAWIO_0_3,requestAWIO_0_2,requestAWIO_0_1,requestAWIO_0_0}; // @[Xbar.scala 64:75]
  assign _T_140 = {requestAWIO_0_12,requestAWIO_0_11,requestAWIO_0_10,requestAWIO_0_9,requestAWIO_0_8,requestAWIO_0_7,requestAWIO_0_6}; // @[Xbar.scala 64:75]
  assign _T_141 = {requestAWIO_0_12,requestAWIO_0_11,requestAWIO_0_10,requestAWIO_0_9,requestAWIO_0_8,requestAWIO_0_7,requestAWIO_0_6,_T_134}; // @[Xbar.scala 64:75]
  assign requestWIO_0_0 = awIn_0_io_deq_bits[0]; // @[Xbar.scala 65:73]
  assign requestWIO_0_1 = awIn_0_io_deq_bits[1]; // @[Xbar.scala 65:73]
  assign requestWIO_0_2 = awIn_0_io_deq_bits[2]; // @[Xbar.scala 65:73]
  assign requestWIO_0_3 = awIn_0_io_deq_bits[3]; // @[Xbar.scala 65:73]
  assign requestWIO_0_4 = awIn_0_io_deq_bits[4]; // @[Xbar.scala 65:73]
  assign requestWIO_0_5 = awIn_0_io_deq_bits[5]; // @[Xbar.scala 65:73]
  assign requestWIO_0_6 = awIn_0_io_deq_bits[6]; // @[Xbar.scala 65:73]
  assign requestWIO_0_7 = awIn_0_io_deq_bits[7]; // @[Xbar.scala 65:73]
  assign requestWIO_0_8 = awIn_0_io_deq_bits[8]; // @[Xbar.scala 65:73]
  assign requestWIO_0_9 = awIn_0_io_deq_bits[9]; // @[Xbar.scala 65:73]
  assign requestWIO_0_10 = awIn_0_io_deq_bits[10]; // @[Xbar.scala 65:73]
  assign requestWIO_0_11 = awIn_0_io_deq_bits[11]; // @[Xbar.scala 65:73]
  assign requestWIO_0_12 = awIn_0_io_deq_bits[12]; // @[Xbar.scala 65:73]
  assign _T_152 = {requestARIO_0_5,requestARIO_0_4,requestARIO_0_3,requestARIO_0_2,requestARIO_0_1,requestARIO_0_0}; // @[Xbar.scala 93:45]
  assign _T_159 = {requestARIO_0_12,requestARIO_0_11,requestARIO_0_10,requestARIO_0_9,requestARIO_0_8,requestARIO_0_7,requestARIO_0_6,_T_152}; // @[Xbar.scala 93:45]
  assign _T_162 = _T_159[12:8] != 5'h0; // @[OneHot.scala 32:14]
  assign _GEN_62 = {{3'd0}, _T_159[12:8]}; // @[OneHot.scala 32:28]
  assign _T_163 = _GEN_62 | _T_159[7:0]; // @[OneHot.scala 32:28]
  assign _T_166 = _T_163[7:4] != 4'h0; // @[OneHot.scala 32:14]
  assign _T_167 = _T_163[7:4] | _T_163[3:0]; // @[OneHot.scala 32:28]
  assign _T_170 = _T_167[3:2] != 2'h0; // @[OneHot.scala 32:14]
  assign _T_171 = _T_167[3:2] | _T_167[1:0]; // @[OneHot.scala 32:28]
  assign _T_175 = {_T_162,_T_166,_T_170,_T_171[1]}; // @[Cat.scala 29:58]
  assign _T_190 = _T_141[12:8] != 5'h0; // @[OneHot.scala 32:14]
  assign _GEN_63 = {{3'd0}, _T_141[12:8]}; // @[OneHot.scala 32:28]
  assign _T_191 = _GEN_63 | _T_141[7:0]; // @[OneHot.scala 32:28]
  assign _T_194 = _T_191[7:4] != 4'h0; // @[OneHot.scala 32:14]
  assign _T_195 = _T_191[7:4] | _T_191[3:0]; // @[OneHot.scala 32:28]
  assign _T_198 = _T_195[3:2] != 2'h0; // @[OneHot.scala 32:14]
  assign _T_199 = _T_195[3:2] | _T_195[1:0]; // @[OneHot.scala 32:28]
  assign _T_203 = {_T_190,_T_194,_T_198,_T_199[1]}; // @[Cat.scala 29:58]
  assign _T_292 = requestARIO_0_0 & auto_out_0_ar_ready; // @[Mux.scala 27:72]
  assign _T_293 = requestARIO_0_1 & auto_out_1_ar_ready; // @[Mux.scala 27:72]
  assign _T_305 = _T_292 | _T_293; // @[Mux.scala 27:72]
  assign _T_294 = requestARIO_0_2 & auto_out_2_ar_ready; // @[Mux.scala 27:72]
  assign _T_306 = _T_305 | _T_294; // @[Mux.scala 27:72]
  assign _T_295 = requestARIO_0_3 & auto_out_3_ar_ready; // @[Mux.scala 27:72]
  assign _T_307 = _T_306 | _T_295; // @[Mux.scala 27:72]
  assign _T_296 = requestARIO_0_4 & auto_out_4_ar_ready; // @[Mux.scala 27:72]
  assign _T_308 = _T_307 | _T_296; // @[Mux.scala 27:72]
  assign _T_297 = requestARIO_0_5 & auto_out_5_ar_ready; // @[Mux.scala 27:72]
  assign _T_309 = _T_308 | _T_297; // @[Mux.scala 27:72]
  assign _T_298 = requestARIO_0_6 & auto_out_6_ar_ready; // @[Mux.scala 27:72]
  assign _T_310 = _T_309 | _T_298; // @[Mux.scala 27:72]
  assign _T_299 = requestARIO_0_7 & auto_out_7_ar_ready; // @[Mux.scala 27:72]
  assign _T_311 = _T_310 | _T_299; // @[Mux.scala 27:72]
  assign _T_300 = requestARIO_0_8 & auto_out_8_ar_ready; // @[Mux.scala 27:72]
  assign _T_312 = _T_311 | _T_300; // @[Mux.scala 27:72]
  assign _T_301 = requestARIO_0_9 & auto_out_9_ar_ready; // @[Mux.scala 27:72]
  assign _T_313 = _T_312 | _T_301; // @[Mux.scala 27:72]
  assign _T_302 = requestARIO_0_10 & auto_out_10_ar_ready; // @[Mux.scala 27:72]
  assign _T_314 = _T_313 | _T_302; // @[Mux.scala 27:72]
  assign _T_303 = requestARIO_0_11 & auto_out_11_ar_ready; // @[Mux.scala 27:72]
  assign _T_315 = _T_314 | _T_303; // @[Mux.scala 27:72]
  assign _T_304 = requestARIO_0_12 & auto_out_12_ar_ready; // @[Mux.scala 27:72]
  assign in_0_ar_ready = _T_315 | _T_304; // @[Mux.scala 27:72]
  assign _T_228 = _T_209 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_227 = _T_210 == _T_175; // @[Xbar.scala 111:75]
  assign _T_229 = _T_228 | _T_227; // @[Xbar.scala 112:34]
  assign _T_230 = _T_209 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_232 = _T_229 & _T_230; // @[Xbar.scala 112:48]
  assign io_in_0_ar_ready = in_0_ar_ready & _T_232; // @[Xbar.scala 130:45]
  assign _T_204 = io_in_0_ar_ready & auto_in_ar_valid; // @[Decoupled.scala 40:37]
  assign _T_399 = auto_out_0_r_valid & requestROI_0_0; // @[Xbar.scala 222:40]
  assign _T_401 = auto_out_1_r_valid & requestROI_1_0; // @[Xbar.scala 222:40]
  assign _T_1023 = _T_399 | _T_401; // @[Xbar.scala 246:36]
  assign _T_403 = auto_out_2_r_valid & requestROI_2_0; // @[Xbar.scala 222:40]
  assign _T_1024 = _T_1023 | _T_403; // @[Xbar.scala 246:36]
  assign _T_405 = auto_out_3_r_valid & requestROI_3_0; // @[Xbar.scala 222:40]
  assign _T_1025 = _T_1024 | _T_405; // @[Xbar.scala 246:36]
  assign _T_407 = auto_out_4_r_valid & requestROI_4_0; // @[Xbar.scala 222:40]
  assign _T_1026 = _T_1025 | _T_407; // @[Xbar.scala 246:36]
  assign _T_409 = auto_out_5_r_valid & requestROI_5_0; // @[Xbar.scala 222:40]
  assign _T_1027 = _T_1026 | _T_409; // @[Xbar.scala 246:36]
  assign _T_411 = auto_out_6_r_valid & requestROI_6_0; // @[Xbar.scala 222:40]
  assign _T_1028 = _T_1027 | _T_411; // @[Xbar.scala 246:36]
  assign _T_413 = auto_out_7_r_valid & requestROI_7_0; // @[Xbar.scala 222:40]
  assign _T_1029 = _T_1028 | _T_413; // @[Xbar.scala 246:36]
  assign _T_415 = auto_out_8_r_valid & requestROI_8_0; // @[Xbar.scala 222:40]
  assign _T_1030 = _T_1029 | _T_415; // @[Xbar.scala 246:36]
  assign _T_417 = auto_out_9_r_valid & requestROI_9_0; // @[Xbar.scala 222:40]
  assign _T_1031 = _T_1030 | _T_417; // @[Xbar.scala 246:36]
  assign _T_419 = auto_out_10_r_valid & requestROI_10_0; // @[Xbar.scala 222:40]
  assign _T_1032 = _T_1031 | _T_419; // @[Xbar.scala 246:36]
  assign _T_421 = auto_out_11_r_valid & requestROI_11_0; // @[Xbar.scala 222:40]
  assign _T_1033 = _T_1032 | _T_421; // @[Xbar.scala 246:36]
  assign _T_423 = auto_out_12_r_valid & requestROI_12_0; // @[Xbar.scala 222:40]
  assign _T_1034 = _T_1033 | _T_423; // @[Xbar.scala 246:36]
  assign _T_1220 = _T_1203_0 & _T_399; // @[Mux.scala 27:72]
  assign _T_1221 = _T_1203_1 & _T_401; // @[Mux.scala 27:72]
  assign _T_1233 = _T_1220 | _T_1221; // @[Mux.scala 27:72]
  assign _T_1222 = _T_1203_2 & _T_403; // @[Mux.scala 27:72]
  assign _T_1234 = _T_1233 | _T_1222; // @[Mux.scala 27:72]
  assign _T_1223 = _T_1203_3 & _T_405; // @[Mux.scala 27:72]
  assign _T_1235 = _T_1234 | _T_1223; // @[Mux.scala 27:72]
  assign _T_1224 = _T_1203_4 & _T_407; // @[Mux.scala 27:72]
  assign _T_1236 = _T_1235 | _T_1224; // @[Mux.scala 27:72]
  assign _T_1225 = _T_1203_5 & _T_409; // @[Mux.scala 27:72]
  assign _T_1237 = _T_1236 | _T_1225; // @[Mux.scala 27:72]
  assign _T_1226 = _T_1203_6 & _T_411; // @[Mux.scala 27:72]
  assign _T_1238 = _T_1237 | _T_1226; // @[Mux.scala 27:72]
  assign _T_1227 = _T_1203_7 & _T_413; // @[Mux.scala 27:72]
  assign _T_1239 = _T_1238 | _T_1227; // @[Mux.scala 27:72]
  assign _T_1228 = _T_1203_8 & _T_415; // @[Mux.scala 27:72]
  assign _T_1240 = _T_1239 | _T_1228; // @[Mux.scala 27:72]
  assign _T_1229 = _T_1203_9 & _T_417; // @[Mux.scala 27:72]
  assign _T_1241 = _T_1240 | _T_1229; // @[Mux.scala 27:72]
  assign _T_1230 = _T_1203_10 & _T_419; // @[Mux.scala 27:72]
  assign _T_1242 = _T_1241 | _T_1230; // @[Mux.scala 27:72]
  assign _T_1231 = _T_1203_11 & _T_421; // @[Mux.scala 27:72]
  assign _T_1243 = _T_1242 | _T_1231; // @[Mux.scala 27:72]
  assign _T_1232 = _T_1203_12 & _T_423; // @[Mux.scala 27:72]
  assign _T_1244 = _T_1243 | _T_1232; // @[Mux.scala 27:72]
  assign in_0_r_valid = _T_1022 ? _T_1034 : _T_1244; // @[Xbar.scala 278:22]
  assign _T_206 = auto_in_r_ready & in_0_r_valid; // @[Decoupled.scala 40:37]
  assign _T_1039 = {_T_409,_T_407,_T_405,_T_403,_T_401,_T_399}; // @[Cat.scala 29:58]
  assign _T_1046 = {_T_423,_T_421,_T_419,_T_417,_T_415,_T_413,_T_411,_T_1039}; // @[Cat.scala 29:58]
  assign _T_1054 = ~_T_1053; // @[Arbiter.scala 21:30]
  assign _T_1055 = _T_1046 & _T_1054; // @[Arbiter.scala 21:28]
  assign _T_1056 = {_T_1055,_T_423,_T_421,_T_419,_T_417,_T_415,_T_413,_T_411,_T_1039}; // @[Cat.scala 29:58]
  assign _GEN_64 = {{1'd0}, _T_1056[25:1]}; // @[package.scala 208:43]
  assign _T_1058 = _T_1056 | _GEN_64; // @[package.scala 208:43]
  assign _GEN_65 = {{2'd0}, _T_1058[25:2]}; // @[package.scala 208:43]
  assign _T_1060 = _T_1058 | _GEN_65; // @[package.scala 208:43]
  assign _GEN_66 = {{4'd0}, _T_1060[25:4]}; // @[package.scala 208:43]
  assign _T_1062 = _T_1060 | _GEN_66; // @[package.scala 208:43]
  assign _GEN_67 = {{8'd0}, _T_1062[25:8]}; // @[package.scala 208:43]
  assign _T_1064 = _T_1062 | _GEN_67; // @[package.scala 208:43]
  assign _T_1067 = {_T_1053, 13'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_68 = {{1'd0}, _T_1064[25:1]}; // @[Arbiter.scala 22:58]
  assign _T_1068 = _GEN_68 | _T_1067; // @[Arbiter.scala 22:58]
  assign _T_1071 = _T_1068[25:13] & _T_1068[12:0]; // @[Arbiter.scala 23:39]
  assign _T_1072 = ~_T_1071; // @[Arbiter.scala 23:18]
  assign _T_1104 = _T_1072[0] & _T_399; // @[Xbar.scala 250:63]
  assign _T_1204_0 = _T_1022 ? _T_1104 : _T_1203_0; // @[Xbar.scala 262:23]
  assign _T_1249 = {auto_out_0_r_bits_id,auto_out_0_r_bits_data,auto_out_0_r_bits_resp,auto_out_0_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1250 = _T_1204_0 ? _T_1249 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1105 = _T_1072[1] & _T_401; // @[Xbar.scala 250:63]
  assign _T_1204_1 = _T_1022 ? _T_1105 : _T_1203_1; // @[Xbar.scala 262:23]
  assign _T_1253 = {auto_out_1_r_bits_id,auto_out_1_r_bits_data,auto_out_1_r_bits_resp,auto_out_1_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1254 = _T_1204_1 ? _T_1253 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1299 = _T_1250 | _T_1254; // @[Mux.scala 27:72]
  assign _T_1106 = _T_1072[2] & _T_403; // @[Xbar.scala 250:63]
  assign _T_1204_2 = _T_1022 ? _T_1106 : _T_1203_2; // @[Xbar.scala 262:23]
  assign _T_1257 = {auto_out_2_r_bits_id,auto_out_2_r_bits_data,auto_out_2_r_bits_resp,auto_out_2_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1258 = _T_1204_2 ? _T_1257 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1300 = _T_1299 | _T_1258; // @[Mux.scala 27:72]
  assign _T_1107 = _T_1072[3] & _T_405; // @[Xbar.scala 250:63]
  assign _T_1204_3 = _T_1022 ? _T_1107 : _T_1203_3; // @[Xbar.scala 262:23]
  assign _T_1261 = {auto_out_3_r_bits_id,auto_out_3_r_bits_data,auto_out_3_r_bits_resp,auto_out_3_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1262 = _T_1204_3 ? _T_1261 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1301 = _T_1300 | _T_1262; // @[Mux.scala 27:72]
  assign _T_1108 = _T_1072[4] & _T_407; // @[Xbar.scala 250:63]
  assign _T_1204_4 = _T_1022 ? _T_1108 : _T_1203_4; // @[Xbar.scala 262:23]
  assign _T_1265 = {auto_out_4_r_bits_id,auto_out_4_r_bits_data,auto_out_4_r_bits_resp,auto_out_4_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1266 = _T_1204_4 ? _T_1265 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1302 = _T_1301 | _T_1266; // @[Mux.scala 27:72]
  assign _T_1109 = _T_1072[5] & _T_409; // @[Xbar.scala 250:63]
  assign _T_1204_5 = _T_1022 ? _T_1109 : _T_1203_5; // @[Xbar.scala 262:23]
  assign _T_1269 = {auto_out_5_r_bits_id,auto_out_5_r_bits_data,auto_out_5_r_bits_resp,auto_out_5_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1270 = _T_1204_5 ? _T_1269 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1303 = _T_1302 | _T_1270; // @[Mux.scala 27:72]
  assign _T_1110 = _T_1072[6] & _T_411; // @[Xbar.scala 250:63]
  assign _T_1204_6 = _T_1022 ? _T_1110 : _T_1203_6; // @[Xbar.scala 262:23]
  assign _T_1273 = {auto_out_6_r_bits_id,auto_out_6_r_bits_data,auto_out_6_r_bits_resp,auto_out_6_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1274 = _T_1204_6 ? _T_1273 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1304 = _T_1303 | _T_1274; // @[Mux.scala 27:72]
  assign _T_1111 = _T_1072[7] & _T_413; // @[Xbar.scala 250:63]
  assign _T_1204_7 = _T_1022 ? _T_1111 : _T_1203_7; // @[Xbar.scala 262:23]
  assign _T_1277 = {auto_out_7_r_bits_id,auto_out_7_r_bits_data,auto_out_7_r_bits_resp,auto_out_7_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1278 = _T_1204_7 ? _T_1277 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1305 = _T_1304 | _T_1278; // @[Mux.scala 27:72]
  assign _T_1112 = _T_1072[8] & _T_415; // @[Xbar.scala 250:63]
  assign _T_1204_8 = _T_1022 ? _T_1112 : _T_1203_8; // @[Xbar.scala 262:23]
  assign _T_1281 = {auto_out_8_r_bits_id,auto_out_8_r_bits_data,auto_out_8_r_bits_resp,auto_out_8_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1282 = _T_1204_8 ? _T_1281 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1306 = _T_1305 | _T_1282; // @[Mux.scala 27:72]
  assign _T_1113 = _T_1072[9] & _T_417; // @[Xbar.scala 250:63]
  assign _T_1204_9 = _T_1022 ? _T_1113 : _T_1203_9; // @[Xbar.scala 262:23]
  assign _T_1285 = {auto_out_9_r_bits_id,auto_out_9_r_bits_data,auto_out_9_r_bits_resp,auto_out_9_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1286 = _T_1204_9 ? _T_1285 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1307 = _T_1306 | _T_1286; // @[Mux.scala 27:72]
  assign _T_1114 = _T_1072[10] & _T_419; // @[Xbar.scala 250:63]
  assign _T_1204_10 = _T_1022 ? _T_1114 : _T_1203_10; // @[Xbar.scala 262:23]
  assign _T_1289 = {auto_out_10_r_bits_id,auto_out_10_r_bits_data,auto_out_10_r_bits_resp,auto_out_10_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1290 = _T_1204_10 ? _T_1289 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1308 = _T_1307 | _T_1290; // @[Mux.scala 27:72]
  assign _T_1115 = _T_1072[11] & _T_421; // @[Xbar.scala 250:63]
  assign _T_1204_11 = _T_1022 ? _T_1115 : _T_1203_11; // @[Xbar.scala 262:23]
  assign _T_1293 = {auto_out_11_r_bits_id,auto_out_11_r_bits_data,auto_out_11_r_bits_resp,auto_out_11_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1294 = _T_1204_11 ? _T_1293 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1309 = _T_1308 | _T_1294; // @[Mux.scala 27:72]
  assign _T_1116 = _T_1072[12] & _T_423; // @[Xbar.scala 250:63]
  assign _T_1204_12 = _T_1022 ? _T_1116 : _T_1203_12; // @[Xbar.scala 262:23]
  assign _T_1297 = {auto_out_12_r_bits_id,auto_out_12_r_bits_data,auto_out_12_r_bits_resp,auto_out_12_r_bits_last}; // @[Mux.scala 27:72]
  assign _T_1298 = _T_1204_12 ? _T_1297 : 36'h0; // @[Mux.scala 27:72]
  assign _T_1310 = _T_1309 | _T_1298; // @[Mux.scala 27:72]
  assign in_0_r_bits_last = _T_1310[0]; // @[Mux.scala 27:72]
  assign _T_208 = _T_206 & in_0_r_bits_last; // @[Xbar.scala 120:45]
  assign _GEN_69 = {{2'd0}, _T_204}; // @[Xbar.scala 106:30]
  assign _T_212 = _T_209 + _GEN_69; // @[Xbar.scala 106:30]
  assign _GEN_70 = {{2'd0}, _T_208}; // @[Xbar.scala 106:48]
  assign _T_214 = _T_212 - _GEN_70; // @[Xbar.scala 106:48]
  assign _T_215 = ~_T_208; // @[Xbar.scala 107:23]
  assign _T_216 = _T_209 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_217 = _T_215 | _T_216; // @[Xbar.scala 107:34]
  assign _T_219 = _T_217 | reset; // @[Xbar.scala 107:22]
  assign _T_220 = ~_T_219; // @[Xbar.scala 107:22]
  assign _T_221 = ~_T_204; // @[Xbar.scala 108:23]
  assign _T_223 = _T_221 | _T_230; // @[Xbar.scala 108:34]
  assign _T_225 = _T_223 | reset; // @[Xbar.scala 108:22]
  assign _T_226 = ~_T_225; // @[Xbar.scala 108:22]
  assign _T_332 = requestAWIO_0_0 & auto_out_0_aw_ready; // @[Mux.scala 27:72]
  assign _T_333 = requestAWIO_0_1 & auto_out_1_aw_ready; // @[Mux.scala 27:72]
  assign _T_345 = _T_332 | _T_333; // @[Mux.scala 27:72]
  assign _T_334 = requestAWIO_0_2 & auto_out_2_aw_ready; // @[Mux.scala 27:72]
  assign _T_346 = _T_345 | _T_334; // @[Mux.scala 27:72]
  assign _T_335 = requestAWIO_0_3 & auto_out_3_aw_ready; // @[Mux.scala 27:72]
  assign _T_347 = _T_346 | _T_335; // @[Mux.scala 27:72]
  assign _T_336 = requestAWIO_0_4 & auto_out_4_aw_ready; // @[Mux.scala 27:72]
  assign _T_348 = _T_347 | _T_336; // @[Mux.scala 27:72]
  assign _T_337 = requestAWIO_0_5 & auto_out_5_aw_ready; // @[Mux.scala 27:72]
  assign _T_349 = _T_348 | _T_337; // @[Mux.scala 27:72]
  assign _T_338 = requestAWIO_0_6 & auto_out_6_aw_ready; // @[Mux.scala 27:72]
  assign _T_350 = _T_349 | _T_338; // @[Mux.scala 27:72]
  assign _T_339 = requestAWIO_0_7 & auto_out_7_aw_ready; // @[Mux.scala 27:72]
  assign _T_351 = _T_350 | _T_339; // @[Mux.scala 27:72]
  assign _T_340 = requestAWIO_0_8 & auto_out_8_aw_ready; // @[Mux.scala 27:72]
  assign _T_352 = _T_351 | _T_340; // @[Mux.scala 27:72]
  assign _T_341 = requestAWIO_0_9 & auto_out_9_aw_ready; // @[Mux.scala 27:72]
  assign _T_353 = _T_352 | _T_341; // @[Mux.scala 27:72]
  assign _T_342 = requestAWIO_0_10 & auto_out_10_aw_ready; // @[Mux.scala 27:72]
  assign _T_354 = _T_353 | _T_342; // @[Mux.scala 27:72]
  assign _T_343 = requestAWIO_0_11 & auto_out_11_aw_ready; // @[Mux.scala 27:72]
  assign _T_355 = _T_354 | _T_343; // @[Mux.scala 27:72]
  assign _T_344 = requestAWIO_0_12 & auto_out_12_aw_ready; // @[Mux.scala 27:72]
  assign in_0_aw_ready = _T_355 | _T_344; // @[Mux.scala 27:72]
  assign _T_267 = _T_263 | awIn_0_io_enq_ready; // @[Xbar.scala 139:57]
  assign _T_268 = in_0_aw_ready & _T_267; // @[Xbar.scala 139:45]
  assign _T_256 = _T_237 == 3'h0; // @[Xbar.scala 112:22]
  assign _T_255 = _T_238 == _T_203; // @[Xbar.scala 111:75]
  assign _T_257 = _T_256 | _T_255; // @[Xbar.scala 112:34]
  assign _T_258 = _T_237 != 3'h7; // @[Xbar.scala 112:80]
  assign _T_260 = _T_257 & _T_258; // @[Xbar.scala 112:48]
  assign io_in_0_aw_ready = _T_268 & _T_260; // @[Xbar.scala 139:82]
  assign _T_233 = io_in_0_aw_ready & auto_in_aw_valid; // @[Decoupled.scala 40:37]
  assign _T_425 = auto_out_0_b_valid & requestBOI_0_0; // @[Xbar.scala 222:40]
  assign _T_427 = auto_out_1_b_valid & requestBOI_1_0; // @[Xbar.scala 222:40]
  assign _T_1318 = _T_425 | _T_427; // @[Xbar.scala 246:36]
  assign _T_429 = auto_out_2_b_valid & requestBOI_2_0; // @[Xbar.scala 222:40]
  assign _T_1319 = _T_1318 | _T_429; // @[Xbar.scala 246:36]
  assign _T_431 = auto_out_3_b_valid & requestBOI_3_0; // @[Xbar.scala 222:40]
  assign _T_1320 = _T_1319 | _T_431; // @[Xbar.scala 246:36]
  assign _T_433 = auto_out_4_b_valid & requestBOI_4_0; // @[Xbar.scala 222:40]
  assign _T_1321 = _T_1320 | _T_433; // @[Xbar.scala 246:36]
  assign _T_435 = auto_out_5_b_valid & requestBOI_5_0; // @[Xbar.scala 222:40]
  assign _T_1322 = _T_1321 | _T_435; // @[Xbar.scala 246:36]
  assign _T_437 = auto_out_6_b_valid & requestBOI_6_0; // @[Xbar.scala 222:40]
  assign _T_1323 = _T_1322 | _T_437; // @[Xbar.scala 246:36]
  assign _T_439 = auto_out_7_b_valid & requestBOI_7_0; // @[Xbar.scala 222:40]
  assign _T_1324 = _T_1323 | _T_439; // @[Xbar.scala 246:36]
  assign _T_441 = auto_out_8_b_valid & requestBOI_8_0; // @[Xbar.scala 222:40]
  assign _T_1325 = _T_1324 | _T_441; // @[Xbar.scala 246:36]
  assign _T_443 = auto_out_9_b_valid & requestBOI_9_0; // @[Xbar.scala 222:40]
  assign _T_1326 = _T_1325 | _T_443; // @[Xbar.scala 246:36]
  assign _T_445 = auto_out_10_b_valid & requestBOI_10_0; // @[Xbar.scala 222:40]
  assign _T_1327 = _T_1326 | _T_445; // @[Xbar.scala 246:36]
  assign _T_447 = auto_out_11_b_valid & requestBOI_11_0; // @[Xbar.scala 222:40]
  assign _T_1328 = _T_1327 | _T_447; // @[Xbar.scala 246:36]
  assign _T_449 = auto_out_12_b_valid & requestBOI_12_0; // @[Xbar.scala 222:40]
  assign _T_1329 = _T_1328 | _T_449; // @[Xbar.scala 246:36]
  assign _T_1515 = _T_1498_0 & _T_425; // @[Mux.scala 27:72]
  assign _T_1516 = _T_1498_1 & _T_427; // @[Mux.scala 27:72]
  assign _T_1528 = _T_1515 | _T_1516; // @[Mux.scala 27:72]
  assign _T_1517 = _T_1498_2 & _T_429; // @[Mux.scala 27:72]
  assign _T_1529 = _T_1528 | _T_1517; // @[Mux.scala 27:72]
  assign _T_1518 = _T_1498_3 & _T_431; // @[Mux.scala 27:72]
  assign _T_1530 = _T_1529 | _T_1518; // @[Mux.scala 27:72]
  assign _T_1519 = _T_1498_4 & _T_433; // @[Mux.scala 27:72]
  assign _T_1531 = _T_1530 | _T_1519; // @[Mux.scala 27:72]
  assign _T_1520 = _T_1498_5 & _T_435; // @[Mux.scala 27:72]
  assign _T_1532 = _T_1531 | _T_1520; // @[Mux.scala 27:72]
  assign _T_1521 = _T_1498_6 & _T_437; // @[Mux.scala 27:72]
  assign _T_1533 = _T_1532 | _T_1521; // @[Mux.scala 27:72]
  assign _T_1522 = _T_1498_7 & _T_439; // @[Mux.scala 27:72]
  assign _T_1534 = _T_1533 | _T_1522; // @[Mux.scala 27:72]
  assign _T_1523 = _T_1498_8 & _T_441; // @[Mux.scala 27:72]
  assign _T_1535 = _T_1534 | _T_1523; // @[Mux.scala 27:72]
  assign _T_1524 = _T_1498_9 & _T_443; // @[Mux.scala 27:72]
  assign _T_1536 = _T_1535 | _T_1524; // @[Mux.scala 27:72]
  assign _T_1525 = _T_1498_10 & _T_445; // @[Mux.scala 27:72]
  assign _T_1537 = _T_1536 | _T_1525; // @[Mux.scala 27:72]
  assign _T_1526 = _T_1498_11 & _T_447; // @[Mux.scala 27:72]
  assign _T_1538 = _T_1537 | _T_1526; // @[Mux.scala 27:72]
  assign _T_1527 = _T_1498_12 & _T_449; // @[Mux.scala 27:72]
  assign _T_1539 = _T_1538 | _T_1527; // @[Mux.scala 27:72]
  assign in_0_b_valid = _T_1317 ? _T_1329 : _T_1539; // @[Xbar.scala 278:22]
  assign _T_235 = auto_in_b_ready & in_0_b_valid; // @[Decoupled.scala 40:37]
  assign _GEN_71 = {{2'd0}, _T_233}; // @[Xbar.scala 106:30]
  assign _T_240 = _T_237 + _GEN_71; // @[Xbar.scala 106:30]
  assign _GEN_72 = {{2'd0}, _T_235}; // @[Xbar.scala 106:48]
  assign _T_242 = _T_240 - _GEN_72; // @[Xbar.scala 106:48]
  assign _T_243 = ~_T_235; // @[Xbar.scala 107:23]
  assign _T_244 = _T_237 != 3'h0; // @[Xbar.scala 107:43]
  assign _T_245 = _T_243 | _T_244; // @[Xbar.scala 107:34]
  assign _T_247 = _T_245 | reset; // @[Xbar.scala 107:22]
  assign _T_248 = ~_T_247; // @[Xbar.scala 107:22]
  assign _T_249 = ~_T_233; // @[Xbar.scala 108:23]
  assign _T_251 = _T_249 | _T_258; // @[Xbar.scala 108:34]
  assign _T_253 = _T_251 | reset; // @[Xbar.scala 108:22]
  assign _T_254 = ~_T_253; // @[Xbar.scala 108:22]
  assign in_0_ar_valid = auto_in_ar_valid & _T_232; // @[Xbar.scala 129:45]
  assign _T_265 = auto_in_aw_valid & _T_267; // @[Xbar.scala 138:45]
  assign in_0_aw_valid = _T_265 & _T_260; // @[Xbar.scala 138:82]
  assign _T_270 = ~_T_263; // @[Xbar.scala 140:54]
  assign _T_272 = awIn_0_io_enq_ready & awIn_0_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_272 | _T_263; // @[Xbar.scala 141:38]
  assign _T_273 = in_0_aw_ready & in_0_aw_valid; // @[Decoupled.scala 40:37]
  assign in_0_w_valid = auto_in_w_valid & awIn_0_io_deq_valid; // @[Xbar.scala 145:43]
  assign _T_372 = requestWIO_0_0 & auto_out_0_w_ready; // @[Mux.scala 27:72]
  assign _T_373 = requestWIO_0_1 & auto_out_1_w_ready; // @[Mux.scala 27:72]
  assign _T_385 = _T_372 | _T_373; // @[Mux.scala 27:72]
  assign _T_374 = requestWIO_0_2 & auto_out_2_w_ready; // @[Mux.scala 27:72]
  assign _T_386 = _T_385 | _T_374; // @[Mux.scala 27:72]
  assign _T_375 = requestWIO_0_3 & auto_out_3_w_ready; // @[Mux.scala 27:72]
  assign _T_387 = _T_386 | _T_375; // @[Mux.scala 27:72]
  assign _T_376 = requestWIO_0_4 & auto_out_4_w_ready; // @[Mux.scala 27:72]
  assign _T_388 = _T_387 | _T_376; // @[Mux.scala 27:72]
  assign _T_377 = requestWIO_0_5 & auto_out_5_w_ready; // @[Mux.scala 27:72]
  assign _T_389 = _T_388 | _T_377; // @[Mux.scala 27:72]
  assign _T_378 = requestWIO_0_6 & auto_out_6_w_ready; // @[Mux.scala 27:72]
  assign _T_390 = _T_389 | _T_378; // @[Mux.scala 27:72]
  assign _T_379 = requestWIO_0_7 & auto_out_7_w_ready; // @[Mux.scala 27:72]
  assign _T_391 = _T_390 | _T_379; // @[Mux.scala 27:72]
  assign _T_380 = requestWIO_0_8 & auto_out_8_w_ready; // @[Mux.scala 27:72]
  assign _T_392 = _T_391 | _T_380; // @[Mux.scala 27:72]
  assign _T_381 = requestWIO_0_9 & auto_out_9_w_ready; // @[Mux.scala 27:72]
  assign _T_393 = _T_392 | _T_381; // @[Mux.scala 27:72]
  assign _T_382 = requestWIO_0_10 & auto_out_10_w_ready; // @[Mux.scala 27:72]
  assign _T_394 = _T_393 | _T_382; // @[Mux.scala 27:72]
  assign _T_383 = requestWIO_0_11 & auto_out_11_w_ready; // @[Mux.scala 27:72]
  assign _T_395 = _T_394 | _T_383; // @[Mux.scala 27:72]
  assign _T_384 = requestWIO_0_12 & auto_out_12_w_ready; // @[Mux.scala 27:72]
  assign in_0_w_ready = _T_395 | _T_384; // @[Mux.scala 27:72]
  assign _T_276 = auto_in_w_valid & auto_in_w_bits_last; // @[Xbar.scala 147:50]
  assign out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[Xbar.scala 222:40]
  assign out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[Xbar.scala 222:40]
  assign out_3_ar_valid = in_0_ar_valid & requestARIO_0_3; // @[Xbar.scala 222:40]
  assign out_4_ar_valid = in_0_ar_valid & requestARIO_0_4; // @[Xbar.scala 222:40]
  assign out_5_ar_valid = in_0_ar_valid & requestARIO_0_5; // @[Xbar.scala 222:40]
  assign out_6_ar_valid = in_0_ar_valid & requestARIO_0_6; // @[Xbar.scala 222:40]
  assign out_7_ar_valid = in_0_ar_valid & requestARIO_0_7; // @[Xbar.scala 222:40]
  assign out_8_ar_valid = in_0_ar_valid & requestARIO_0_8; // @[Xbar.scala 222:40]
  assign out_9_ar_valid = in_0_ar_valid & requestARIO_0_9; // @[Xbar.scala 222:40]
  assign out_10_ar_valid = in_0_ar_valid & requestARIO_0_10; // @[Xbar.scala 222:40]
  assign out_11_ar_valid = in_0_ar_valid & requestARIO_0_11; // @[Xbar.scala 222:40]
  assign out_12_ar_valid = in_0_ar_valid & requestARIO_0_12; // @[Xbar.scala 222:40]
  assign out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[Xbar.scala 222:40]
  assign out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[Xbar.scala 222:40]
  assign out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[Xbar.scala 222:40]
  assign out_3_aw_valid = in_0_aw_valid & requestAWIO_0_3; // @[Xbar.scala 222:40]
  assign out_4_aw_valid = in_0_aw_valid & requestAWIO_0_4; // @[Xbar.scala 222:40]
  assign out_5_aw_valid = in_0_aw_valid & requestAWIO_0_5; // @[Xbar.scala 222:40]
  assign out_6_aw_valid = in_0_aw_valid & requestAWIO_0_6; // @[Xbar.scala 222:40]
  assign out_7_aw_valid = in_0_aw_valid & requestAWIO_0_7; // @[Xbar.scala 222:40]
  assign out_8_aw_valid = in_0_aw_valid & requestAWIO_0_8; // @[Xbar.scala 222:40]
  assign out_9_aw_valid = in_0_aw_valid & requestAWIO_0_9; // @[Xbar.scala 222:40]
  assign out_10_aw_valid = in_0_aw_valid & requestAWIO_0_10; // @[Xbar.scala 222:40]
  assign out_11_aw_valid = in_0_aw_valid & requestAWIO_0_11; // @[Xbar.scala 222:40]
  assign out_12_aw_valid = in_0_aw_valid & requestAWIO_0_12; // @[Xbar.scala 222:40]
  assign _T_456 = ~out_0_aw_valid; // @[Xbar.scala 256:60]
  assign _T_462 = _T_456 | out_0_aw_valid; // @[Xbar.scala 258:23]
  assign _T_464 = _T_462 | reset; // @[Xbar.scala 258:12]
  assign _T_465 = ~_T_464; // @[Xbar.scala 258:12]
  assign _T_477 = ~out_0_ar_valid; // @[Xbar.scala 256:60]
  assign _T_483 = _T_477 | out_0_ar_valid; // @[Xbar.scala 258:23]
  assign _T_485 = _T_483 | reset; // @[Xbar.scala 258:12]
  assign _T_486 = ~_T_485; // @[Xbar.scala 258:12]
  assign _T_500 = ~out_1_aw_valid; // @[Xbar.scala 256:60]
  assign _T_506 = _T_500 | out_1_aw_valid; // @[Xbar.scala 258:23]
  assign _T_508 = _T_506 | reset; // @[Xbar.scala 258:12]
  assign _T_509 = ~_T_508; // @[Xbar.scala 258:12]
  assign _T_521 = ~out_1_ar_valid; // @[Xbar.scala 256:60]
  assign _T_527 = _T_521 | out_1_ar_valid; // @[Xbar.scala 258:23]
  assign _T_529 = _T_527 | reset; // @[Xbar.scala 258:12]
  assign _T_530 = ~_T_529; // @[Xbar.scala 258:12]
  assign _T_544 = ~out_2_aw_valid; // @[Xbar.scala 256:60]
  assign _T_550 = _T_544 | out_2_aw_valid; // @[Xbar.scala 258:23]
  assign _T_552 = _T_550 | reset; // @[Xbar.scala 258:12]
  assign _T_553 = ~_T_552; // @[Xbar.scala 258:12]
  assign _T_565 = ~out_2_ar_valid; // @[Xbar.scala 256:60]
  assign _T_571 = _T_565 | out_2_ar_valid; // @[Xbar.scala 258:23]
  assign _T_573 = _T_571 | reset; // @[Xbar.scala 258:12]
  assign _T_574 = ~_T_573; // @[Xbar.scala 258:12]
  assign _T_588 = ~out_3_aw_valid; // @[Xbar.scala 256:60]
  assign _T_594 = _T_588 | out_3_aw_valid; // @[Xbar.scala 258:23]
  assign _T_596 = _T_594 | reset; // @[Xbar.scala 258:12]
  assign _T_597 = ~_T_596; // @[Xbar.scala 258:12]
  assign _T_609 = ~out_3_ar_valid; // @[Xbar.scala 256:60]
  assign _T_615 = _T_609 | out_3_ar_valid; // @[Xbar.scala 258:23]
  assign _T_617 = _T_615 | reset; // @[Xbar.scala 258:12]
  assign _T_618 = ~_T_617; // @[Xbar.scala 258:12]
  assign _T_632 = ~out_4_aw_valid; // @[Xbar.scala 256:60]
  assign _T_638 = _T_632 | out_4_aw_valid; // @[Xbar.scala 258:23]
  assign _T_640 = _T_638 | reset; // @[Xbar.scala 258:12]
  assign _T_641 = ~_T_640; // @[Xbar.scala 258:12]
  assign _T_653 = ~out_4_ar_valid; // @[Xbar.scala 256:60]
  assign _T_659 = _T_653 | out_4_ar_valid; // @[Xbar.scala 258:23]
  assign _T_661 = _T_659 | reset; // @[Xbar.scala 258:12]
  assign _T_662 = ~_T_661; // @[Xbar.scala 258:12]
  assign _T_676 = ~out_5_aw_valid; // @[Xbar.scala 256:60]
  assign _T_682 = _T_676 | out_5_aw_valid; // @[Xbar.scala 258:23]
  assign _T_684 = _T_682 | reset; // @[Xbar.scala 258:12]
  assign _T_685 = ~_T_684; // @[Xbar.scala 258:12]
  assign _T_697 = ~out_5_ar_valid; // @[Xbar.scala 256:60]
  assign _T_703 = _T_697 | out_5_ar_valid; // @[Xbar.scala 258:23]
  assign _T_705 = _T_703 | reset; // @[Xbar.scala 258:12]
  assign _T_706 = ~_T_705; // @[Xbar.scala 258:12]
  assign _T_720 = ~out_6_aw_valid; // @[Xbar.scala 256:60]
  assign _T_726 = _T_720 | out_6_aw_valid; // @[Xbar.scala 258:23]
  assign _T_728 = _T_726 | reset; // @[Xbar.scala 258:12]
  assign _T_729 = ~_T_728; // @[Xbar.scala 258:12]
  assign _T_741 = ~out_6_ar_valid; // @[Xbar.scala 256:60]
  assign _T_747 = _T_741 | out_6_ar_valid; // @[Xbar.scala 258:23]
  assign _T_749 = _T_747 | reset; // @[Xbar.scala 258:12]
  assign _T_750 = ~_T_749; // @[Xbar.scala 258:12]
  assign _T_764 = ~out_7_aw_valid; // @[Xbar.scala 256:60]
  assign _T_770 = _T_764 | out_7_aw_valid; // @[Xbar.scala 258:23]
  assign _T_772 = _T_770 | reset; // @[Xbar.scala 258:12]
  assign _T_773 = ~_T_772; // @[Xbar.scala 258:12]
  assign _T_785 = ~out_7_ar_valid; // @[Xbar.scala 256:60]
  assign _T_791 = _T_785 | out_7_ar_valid; // @[Xbar.scala 258:23]
  assign _T_793 = _T_791 | reset; // @[Xbar.scala 258:12]
  assign _T_794 = ~_T_793; // @[Xbar.scala 258:12]
  assign _T_808 = ~out_8_aw_valid; // @[Xbar.scala 256:60]
  assign _T_814 = _T_808 | out_8_aw_valid; // @[Xbar.scala 258:23]
  assign _T_816 = _T_814 | reset; // @[Xbar.scala 258:12]
  assign _T_817 = ~_T_816; // @[Xbar.scala 258:12]
  assign _T_829 = ~out_8_ar_valid; // @[Xbar.scala 256:60]
  assign _T_835 = _T_829 | out_8_ar_valid; // @[Xbar.scala 258:23]
  assign _T_837 = _T_835 | reset; // @[Xbar.scala 258:12]
  assign _T_838 = ~_T_837; // @[Xbar.scala 258:12]
  assign _T_852 = ~out_9_aw_valid; // @[Xbar.scala 256:60]
  assign _T_858 = _T_852 | out_9_aw_valid; // @[Xbar.scala 258:23]
  assign _T_860 = _T_858 | reset; // @[Xbar.scala 258:12]
  assign _T_861 = ~_T_860; // @[Xbar.scala 258:12]
  assign _T_873 = ~out_9_ar_valid; // @[Xbar.scala 256:60]
  assign _T_879 = _T_873 | out_9_ar_valid; // @[Xbar.scala 258:23]
  assign _T_881 = _T_879 | reset; // @[Xbar.scala 258:12]
  assign _T_882 = ~_T_881; // @[Xbar.scala 258:12]
  assign _T_896 = ~out_10_aw_valid; // @[Xbar.scala 256:60]
  assign _T_902 = _T_896 | out_10_aw_valid; // @[Xbar.scala 258:23]
  assign _T_904 = _T_902 | reset; // @[Xbar.scala 258:12]
  assign _T_905 = ~_T_904; // @[Xbar.scala 258:12]
  assign _T_917 = ~out_10_ar_valid; // @[Xbar.scala 256:60]
  assign _T_923 = _T_917 | out_10_ar_valid; // @[Xbar.scala 258:23]
  assign _T_925 = _T_923 | reset; // @[Xbar.scala 258:12]
  assign _T_926 = ~_T_925; // @[Xbar.scala 258:12]
  assign _T_940 = ~out_11_aw_valid; // @[Xbar.scala 256:60]
  assign _T_946 = _T_940 | out_11_aw_valid; // @[Xbar.scala 258:23]
  assign _T_948 = _T_946 | reset; // @[Xbar.scala 258:12]
  assign _T_949 = ~_T_948; // @[Xbar.scala 258:12]
  assign _T_961 = ~out_11_ar_valid; // @[Xbar.scala 256:60]
  assign _T_967 = _T_961 | out_11_ar_valid; // @[Xbar.scala 258:23]
  assign _T_969 = _T_967 | reset; // @[Xbar.scala 258:12]
  assign _T_970 = ~_T_969; // @[Xbar.scala 258:12]
  assign _T_984 = ~out_12_aw_valid; // @[Xbar.scala 256:60]
  assign _T_990 = _T_984 | out_12_aw_valid; // @[Xbar.scala 258:23]
  assign _T_992 = _T_990 | reset; // @[Xbar.scala 258:12]
  assign _T_993 = ~_T_992; // @[Xbar.scala 258:12]
  assign _T_1005 = ~out_12_ar_valid; // @[Xbar.scala 256:60]
  assign _T_1011 = _T_1005 | out_12_ar_valid; // @[Xbar.scala 258:23]
  assign _T_1013 = _T_1011 | reset; // @[Xbar.scala 258:12]
  assign _T_1014 = ~_T_1013; // @[Xbar.scala 258:12]
  assign _T_1073 = _T_1046 != 13'h0; // @[Arbiter.scala 24:27]
  assign _T_1074 = _T_1022 & _T_1073; // @[Arbiter.scala 24:18]
  assign _T_1075 = _T_1072 & _T_1046; // @[Arbiter.scala 25:29]
  assign _T_1076 = {_T_1075, 1'h0}; // @[package.scala 199:48]
  assign _T_1078 = _T_1075 | _T_1076[12:0]; // @[package.scala 199:43]
  assign _T_1079 = {_T_1078, 2'h0}; // @[package.scala 199:48]
  assign _T_1081 = _T_1078 | _T_1079[12:0]; // @[package.scala 199:43]
  assign _T_1082 = {_T_1081, 4'h0}; // @[package.scala 199:48]
  assign _T_1084 = _T_1081 | _T_1082[12:0]; // @[package.scala 199:43]
  assign _T_1085 = {_T_1084, 8'h0}; // @[package.scala 199:48]
  assign _T_1087 = _T_1084 | _T_1085[12:0]; // @[package.scala 199:43]
  assign _T_1119 = _T_1104 | _T_1105; // @[Xbar.scala 255:50]
  assign _T_1120 = _T_1119 | _T_1106; // @[Xbar.scala 255:50]
  assign _T_1121 = _T_1120 | _T_1107; // @[Xbar.scala 255:50]
  assign _T_1122 = _T_1121 | _T_1108; // @[Xbar.scala 255:50]
  assign _T_1123 = _T_1122 | _T_1109; // @[Xbar.scala 255:50]
  assign _T_1124 = _T_1123 | _T_1110; // @[Xbar.scala 255:50]
  assign _T_1125 = _T_1124 | _T_1111; // @[Xbar.scala 255:50]
  assign _T_1126 = _T_1125 | _T_1112; // @[Xbar.scala 255:50]
  assign _T_1127 = _T_1126 | _T_1113; // @[Xbar.scala 255:50]
  assign _T_1128 = _T_1127 | _T_1114; // @[Xbar.scala 255:50]
  assign _T_1129 = _T_1128 | _T_1115; // @[Xbar.scala 255:50]
  assign _T_1130 = _T_1129 | _T_1116; // @[Xbar.scala 255:50]
  assign _T_1132 = ~_T_1104; // @[Xbar.scala 256:60]
  assign _T_1135 = ~_T_1105; // @[Xbar.scala 256:60]
  assign _T_1136 = _T_1132 | _T_1135; // @[Xbar.scala 256:57]
  assign _T_1137 = ~_T_1119; // @[Xbar.scala 256:54]
  assign _T_1138 = ~_T_1106; // @[Xbar.scala 256:60]
  assign _T_1139 = _T_1137 | _T_1138; // @[Xbar.scala 256:57]
  assign _T_1140 = ~_T_1120; // @[Xbar.scala 256:54]
  assign _T_1141 = ~_T_1107; // @[Xbar.scala 256:60]
  assign _T_1142 = _T_1140 | _T_1141; // @[Xbar.scala 256:57]
  assign _T_1143 = ~_T_1121; // @[Xbar.scala 256:54]
  assign _T_1144 = ~_T_1108; // @[Xbar.scala 256:60]
  assign _T_1145 = _T_1143 | _T_1144; // @[Xbar.scala 256:57]
  assign _T_1146 = ~_T_1122; // @[Xbar.scala 256:54]
  assign _T_1147 = ~_T_1109; // @[Xbar.scala 256:60]
  assign _T_1148 = _T_1146 | _T_1147; // @[Xbar.scala 256:57]
  assign _T_1149 = ~_T_1123; // @[Xbar.scala 256:54]
  assign _T_1150 = ~_T_1110; // @[Xbar.scala 256:60]
  assign _T_1151 = _T_1149 | _T_1150; // @[Xbar.scala 256:57]
  assign _T_1152 = ~_T_1124; // @[Xbar.scala 256:54]
  assign _T_1153 = ~_T_1111; // @[Xbar.scala 256:60]
  assign _T_1154 = _T_1152 | _T_1153; // @[Xbar.scala 256:57]
  assign _T_1155 = ~_T_1125; // @[Xbar.scala 256:54]
  assign _T_1156 = ~_T_1112; // @[Xbar.scala 256:60]
  assign _T_1157 = _T_1155 | _T_1156; // @[Xbar.scala 256:57]
  assign _T_1158 = ~_T_1126; // @[Xbar.scala 256:54]
  assign _T_1159 = ~_T_1113; // @[Xbar.scala 256:60]
  assign _T_1160 = _T_1158 | _T_1159; // @[Xbar.scala 256:57]
  assign _T_1161 = ~_T_1127; // @[Xbar.scala 256:54]
  assign _T_1162 = ~_T_1114; // @[Xbar.scala 256:60]
  assign _T_1163 = _T_1161 | _T_1162; // @[Xbar.scala 256:57]
  assign _T_1164 = ~_T_1128; // @[Xbar.scala 256:54]
  assign _T_1165 = ~_T_1115; // @[Xbar.scala 256:60]
  assign _T_1166 = _T_1164 | _T_1165; // @[Xbar.scala 256:57]
  assign _T_1167 = ~_T_1129; // @[Xbar.scala 256:54]
  assign _T_1168 = ~_T_1116; // @[Xbar.scala 256:60]
  assign _T_1169 = _T_1167 | _T_1168; // @[Xbar.scala 256:57]
  assign _T_1171 = _T_1136 & _T_1139; // @[Xbar.scala 256:75]
  assign _T_1172 = _T_1171 & _T_1142; // @[Xbar.scala 256:75]
  assign _T_1173 = _T_1172 & _T_1145; // @[Xbar.scala 256:75]
  assign _T_1174 = _T_1173 & _T_1148; // @[Xbar.scala 256:75]
  assign _T_1175 = _T_1174 & _T_1151; // @[Xbar.scala 256:75]
  assign _T_1176 = _T_1175 & _T_1154; // @[Xbar.scala 256:75]
  assign _T_1177 = _T_1176 & _T_1157; // @[Xbar.scala 256:75]
  assign _T_1178 = _T_1177 & _T_1160; // @[Xbar.scala 256:75]
  assign _T_1179 = _T_1178 & _T_1163; // @[Xbar.scala 256:75]
  assign _T_1180 = _T_1179 & _T_1166; // @[Xbar.scala 256:75]
  assign _T_1181 = _T_1180 & _T_1169; // @[Xbar.scala 256:75]
  assign _T_1183 = _T_1181 | reset; // @[Xbar.scala 256:11]
  assign _T_1184 = ~_T_1183; // @[Xbar.scala 256:11]
  assign _T_1185 = ~_T_1034; // @[Xbar.scala 258:13]
  assign _T_1198 = _T_1185 | _T_1130; // @[Xbar.scala 258:23]
  assign _T_1200 = _T_1198 | reset; // @[Xbar.scala 258:12]
  assign _T_1201 = ~_T_1200; // @[Xbar.scala 258:12]
  assign _GEN_57 = _T_1034 ? 1'h0 : _T_1022; // @[Xbar.scala 266:21]
  assign _GEN_58 = _T_206 | _GEN_57; // @[Xbar.scala 267:24]
  assign _T_1206_0 = _T_1022 ? _T_1072[0] : _T_1203_0; // @[Xbar.scala 270:24]
  assign _T_1206_1 = _T_1022 ? _T_1072[1] : _T_1203_1; // @[Xbar.scala 270:24]
  assign _T_1206_2 = _T_1022 ? _T_1072[2] : _T_1203_2; // @[Xbar.scala 270:24]
  assign _T_1206_3 = _T_1022 ? _T_1072[3] : _T_1203_3; // @[Xbar.scala 270:24]
  assign _T_1206_4 = _T_1022 ? _T_1072[4] : _T_1203_4; // @[Xbar.scala 270:24]
  assign _T_1206_5 = _T_1022 ? _T_1072[5] : _T_1203_5; // @[Xbar.scala 270:24]
  assign _T_1206_6 = _T_1022 ? _T_1072[6] : _T_1203_6; // @[Xbar.scala 270:24]
  assign _T_1206_7 = _T_1022 ? _T_1072[7] : _T_1203_7; // @[Xbar.scala 270:24]
  assign _T_1206_8 = _T_1022 ? _T_1072[8] : _T_1203_8; // @[Xbar.scala 270:24]
  assign _T_1206_9 = _T_1022 ? _T_1072[9] : _T_1203_9; // @[Xbar.scala 270:24]
  assign _T_1206_10 = _T_1022 ? _T_1072[10] : _T_1203_10; // @[Xbar.scala 270:24]
  assign _T_1206_11 = _T_1022 ? _T_1072[11] : _T_1203_11; // @[Xbar.scala 270:24]
  assign _T_1206_12 = _T_1022 ? _T_1072[12] : _T_1203_12; // @[Xbar.scala 270:24]
  assign _T_1334 = {_T_435,_T_433,_T_431,_T_429,_T_427,_T_425}; // @[Cat.scala 29:58]
  assign _T_1341 = {_T_449,_T_447,_T_445,_T_443,_T_441,_T_439,_T_437,_T_1334}; // @[Cat.scala 29:58]
  assign _T_1349 = ~_T_1348; // @[Arbiter.scala 21:30]
  assign _T_1350 = _T_1341 & _T_1349; // @[Arbiter.scala 21:28]
  assign _T_1351 = {_T_1350,_T_449,_T_447,_T_445,_T_443,_T_441,_T_439,_T_437,_T_1334}; // @[Cat.scala 29:58]
  assign _GEN_73 = {{1'd0}, _T_1351[25:1]}; // @[package.scala 208:43]
  assign _T_1353 = _T_1351 | _GEN_73; // @[package.scala 208:43]
  assign _GEN_74 = {{2'd0}, _T_1353[25:2]}; // @[package.scala 208:43]
  assign _T_1355 = _T_1353 | _GEN_74; // @[package.scala 208:43]
  assign _GEN_75 = {{4'd0}, _T_1355[25:4]}; // @[package.scala 208:43]
  assign _T_1357 = _T_1355 | _GEN_75; // @[package.scala 208:43]
  assign _GEN_76 = {{8'd0}, _T_1357[25:8]}; // @[package.scala 208:43]
  assign _T_1359 = _T_1357 | _GEN_76; // @[package.scala 208:43]
  assign _T_1362 = {_T_1348, 13'h0}; // @[Arbiter.scala 22:66]
  assign _GEN_77 = {{1'd0}, _T_1359[25:1]}; // @[Arbiter.scala 22:58]
  assign _T_1363 = _GEN_77 | _T_1362; // @[Arbiter.scala 22:58]
  assign _T_1366 = _T_1363[25:13] & _T_1363[12:0]; // @[Arbiter.scala 23:39]
  assign _T_1367 = ~_T_1366; // @[Arbiter.scala 23:18]
  assign _T_1368 = _T_1341 != 13'h0; // @[Arbiter.scala 24:27]
  assign _T_1369 = _T_1317 & _T_1368; // @[Arbiter.scala 24:18]
  assign _T_1370 = _T_1367 & _T_1341; // @[Arbiter.scala 25:29]
  assign _T_1371 = {_T_1370, 1'h0}; // @[package.scala 199:48]
  assign _T_1373 = _T_1370 | _T_1371[12:0]; // @[package.scala 199:43]
  assign _T_1374 = {_T_1373, 2'h0}; // @[package.scala 199:48]
  assign _T_1376 = _T_1373 | _T_1374[12:0]; // @[package.scala 199:43]
  assign _T_1377 = {_T_1376, 4'h0}; // @[package.scala 199:48]
  assign _T_1379 = _T_1376 | _T_1377[12:0]; // @[package.scala 199:43]
  assign _T_1380 = {_T_1379, 8'h0}; // @[package.scala 199:48]
  assign _T_1382 = _T_1379 | _T_1380[12:0]; // @[package.scala 199:43]
  assign _T_1399 = _T_1367[0] & _T_425; // @[Xbar.scala 250:63]
  assign _T_1400 = _T_1367[1] & _T_427; // @[Xbar.scala 250:63]
  assign _T_1401 = _T_1367[2] & _T_429; // @[Xbar.scala 250:63]
  assign _T_1402 = _T_1367[3] & _T_431; // @[Xbar.scala 250:63]
  assign _T_1403 = _T_1367[4] & _T_433; // @[Xbar.scala 250:63]
  assign _T_1404 = _T_1367[5] & _T_435; // @[Xbar.scala 250:63]
  assign _T_1405 = _T_1367[6] & _T_437; // @[Xbar.scala 250:63]
  assign _T_1406 = _T_1367[7] & _T_439; // @[Xbar.scala 250:63]
  assign _T_1407 = _T_1367[8] & _T_441; // @[Xbar.scala 250:63]
  assign _T_1408 = _T_1367[9] & _T_443; // @[Xbar.scala 250:63]
  assign _T_1409 = _T_1367[10] & _T_445; // @[Xbar.scala 250:63]
  assign _T_1410 = _T_1367[11] & _T_447; // @[Xbar.scala 250:63]
  assign _T_1411 = _T_1367[12] & _T_449; // @[Xbar.scala 250:63]
  assign _T_1414 = _T_1399 | _T_1400; // @[Xbar.scala 255:50]
  assign _T_1415 = _T_1414 | _T_1401; // @[Xbar.scala 255:50]
  assign _T_1416 = _T_1415 | _T_1402; // @[Xbar.scala 255:50]
  assign _T_1417 = _T_1416 | _T_1403; // @[Xbar.scala 255:50]
  assign _T_1418 = _T_1417 | _T_1404; // @[Xbar.scala 255:50]
  assign _T_1419 = _T_1418 | _T_1405; // @[Xbar.scala 255:50]
  assign _T_1420 = _T_1419 | _T_1406; // @[Xbar.scala 255:50]
  assign _T_1421 = _T_1420 | _T_1407; // @[Xbar.scala 255:50]
  assign _T_1422 = _T_1421 | _T_1408; // @[Xbar.scala 255:50]
  assign _T_1423 = _T_1422 | _T_1409; // @[Xbar.scala 255:50]
  assign _T_1424 = _T_1423 | _T_1410; // @[Xbar.scala 255:50]
  assign _T_1425 = _T_1424 | _T_1411; // @[Xbar.scala 255:50]
  assign _T_1427 = ~_T_1399; // @[Xbar.scala 256:60]
  assign _T_1430 = ~_T_1400; // @[Xbar.scala 256:60]
  assign _T_1431 = _T_1427 | _T_1430; // @[Xbar.scala 256:57]
  assign _T_1432 = ~_T_1414; // @[Xbar.scala 256:54]
  assign _T_1433 = ~_T_1401; // @[Xbar.scala 256:60]
  assign _T_1434 = _T_1432 | _T_1433; // @[Xbar.scala 256:57]
  assign _T_1435 = ~_T_1415; // @[Xbar.scala 256:54]
  assign _T_1436 = ~_T_1402; // @[Xbar.scala 256:60]
  assign _T_1437 = _T_1435 | _T_1436; // @[Xbar.scala 256:57]
  assign _T_1438 = ~_T_1416; // @[Xbar.scala 256:54]
  assign _T_1439 = ~_T_1403; // @[Xbar.scala 256:60]
  assign _T_1440 = _T_1438 | _T_1439; // @[Xbar.scala 256:57]
  assign _T_1441 = ~_T_1417; // @[Xbar.scala 256:54]
  assign _T_1442 = ~_T_1404; // @[Xbar.scala 256:60]
  assign _T_1443 = _T_1441 | _T_1442; // @[Xbar.scala 256:57]
  assign _T_1444 = ~_T_1418; // @[Xbar.scala 256:54]
  assign _T_1445 = ~_T_1405; // @[Xbar.scala 256:60]
  assign _T_1446 = _T_1444 | _T_1445; // @[Xbar.scala 256:57]
  assign _T_1447 = ~_T_1419; // @[Xbar.scala 256:54]
  assign _T_1448 = ~_T_1406; // @[Xbar.scala 256:60]
  assign _T_1449 = _T_1447 | _T_1448; // @[Xbar.scala 256:57]
  assign _T_1450 = ~_T_1420; // @[Xbar.scala 256:54]
  assign _T_1451 = ~_T_1407; // @[Xbar.scala 256:60]
  assign _T_1452 = _T_1450 | _T_1451; // @[Xbar.scala 256:57]
  assign _T_1453 = ~_T_1421; // @[Xbar.scala 256:54]
  assign _T_1454 = ~_T_1408; // @[Xbar.scala 256:60]
  assign _T_1455 = _T_1453 | _T_1454; // @[Xbar.scala 256:57]
  assign _T_1456 = ~_T_1422; // @[Xbar.scala 256:54]
  assign _T_1457 = ~_T_1409; // @[Xbar.scala 256:60]
  assign _T_1458 = _T_1456 | _T_1457; // @[Xbar.scala 256:57]
  assign _T_1459 = ~_T_1423; // @[Xbar.scala 256:54]
  assign _T_1460 = ~_T_1410; // @[Xbar.scala 256:60]
  assign _T_1461 = _T_1459 | _T_1460; // @[Xbar.scala 256:57]
  assign _T_1462 = ~_T_1424; // @[Xbar.scala 256:54]
  assign _T_1463 = ~_T_1411; // @[Xbar.scala 256:60]
  assign _T_1464 = _T_1462 | _T_1463; // @[Xbar.scala 256:57]
  assign _T_1466 = _T_1431 & _T_1434; // @[Xbar.scala 256:75]
  assign _T_1467 = _T_1466 & _T_1437; // @[Xbar.scala 256:75]
  assign _T_1468 = _T_1467 & _T_1440; // @[Xbar.scala 256:75]
  assign _T_1469 = _T_1468 & _T_1443; // @[Xbar.scala 256:75]
  assign _T_1470 = _T_1469 & _T_1446; // @[Xbar.scala 256:75]
  assign _T_1471 = _T_1470 & _T_1449; // @[Xbar.scala 256:75]
  assign _T_1472 = _T_1471 & _T_1452; // @[Xbar.scala 256:75]
  assign _T_1473 = _T_1472 & _T_1455; // @[Xbar.scala 256:75]
  assign _T_1474 = _T_1473 & _T_1458; // @[Xbar.scala 256:75]
  assign _T_1475 = _T_1474 & _T_1461; // @[Xbar.scala 256:75]
  assign _T_1476 = _T_1475 & _T_1464; // @[Xbar.scala 256:75]
  assign _T_1478 = _T_1476 | reset; // @[Xbar.scala 256:11]
  assign _T_1479 = ~_T_1478; // @[Xbar.scala 256:11]
  assign _T_1480 = ~_T_1329; // @[Xbar.scala 258:13]
  assign _T_1493 = _T_1480 | _T_1425; // @[Xbar.scala 258:23]
  assign _T_1495 = _T_1493 | reset; // @[Xbar.scala 258:12]
  assign _T_1496 = ~_T_1495; // @[Xbar.scala 258:12]
  assign _T_1499_0 = _T_1317 ? _T_1399 : _T_1498_0; // @[Xbar.scala 262:23]
  assign _T_1499_1 = _T_1317 ? _T_1400 : _T_1498_1; // @[Xbar.scala 262:23]
  assign _T_1499_2 = _T_1317 ? _T_1401 : _T_1498_2; // @[Xbar.scala 262:23]
  assign _T_1499_3 = _T_1317 ? _T_1402 : _T_1498_3; // @[Xbar.scala 262:23]
  assign _T_1499_4 = _T_1317 ? _T_1403 : _T_1498_4; // @[Xbar.scala 262:23]
  assign _T_1499_5 = _T_1317 ? _T_1404 : _T_1498_5; // @[Xbar.scala 262:23]
  assign _T_1499_6 = _T_1317 ? _T_1405 : _T_1498_6; // @[Xbar.scala 262:23]
  assign _T_1499_7 = _T_1317 ? _T_1406 : _T_1498_7; // @[Xbar.scala 262:23]
  assign _T_1499_8 = _T_1317 ? _T_1407 : _T_1498_8; // @[Xbar.scala 262:23]
  assign _T_1499_9 = _T_1317 ? _T_1408 : _T_1498_9; // @[Xbar.scala 262:23]
  assign _T_1499_10 = _T_1317 ? _T_1409 : _T_1498_10; // @[Xbar.scala 262:23]
  assign _T_1499_11 = _T_1317 ? _T_1410 : _T_1498_11; // @[Xbar.scala 262:23]
  assign _T_1499_12 = _T_1317 ? _T_1411 : _T_1498_12; // @[Xbar.scala 262:23]
  assign _GEN_60 = _T_1329 ? 1'h0 : _T_1317; // @[Xbar.scala 266:21]
  assign _GEN_61 = _T_235 | _GEN_60; // @[Xbar.scala 267:24]
  assign _T_1501_0 = _T_1317 ? _T_1367[0] : _T_1498_0; // @[Xbar.scala 270:24]
  assign _T_1501_1 = _T_1317 ? _T_1367[1] : _T_1498_1; // @[Xbar.scala 270:24]
  assign _T_1501_2 = _T_1317 ? _T_1367[2] : _T_1498_2; // @[Xbar.scala 270:24]
  assign _T_1501_3 = _T_1317 ? _T_1367[3] : _T_1498_3; // @[Xbar.scala 270:24]
  assign _T_1501_4 = _T_1317 ? _T_1367[4] : _T_1498_4; // @[Xbar.scala 270:24]
  assign _T_1501_5 = _T_1317 ? _T_1367[5] : _T_1498_5; // @[Xbar.scala 270:24]
  assign _T_1501_6 = _T_1317 ? _T_1367[6] : _T_1498_6; // @[Xbar.scala 270:24]
  assign _T_1501_7 = _T_1317 ? _T_1367[7] : _T_1498_7; // @[Xbar.scala 270:24]
  assign _T_1501_8 = _T_1317 ? _T_1367[8] : _T_1498_8; // @[Xbar.scala 270:24]
  assign _T_1501_9 = _T_1317 ? _T_1367[9] : _T_1498_9; // @[Xbar.scala 270:24]
  assign _T_1501_10 = _T_1317 ? _T_1367[10] : _T_1498_10; // @[Xbar.scala 270:24]
  assign _T_1501_11 = _T_1317 ? _T_1367[11] : _T_1498_11; // @[Xbar.scala 270:24]
  assign _T_1501_12 = _T_1317 ? _T_1367[12] : _T_1498_12; // @[Xbar.scala 270:24]
  assign _T_1542 = {auto_out_0_b_bits_id,auto_out_0_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1543 = _T_1499_0 ? _T_1542 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1544 = {auto_out_1_b_bits_id,auto_out_1_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1545 = _T_1499_1 ? _T_1544 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1546 = {auto_out_2_b_bits_id,auto_out_2_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1547 = _T_1499_2 ? _T_1546 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1548 = {auto_out_3_b_bits_id,auto_out_3_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1549 = _T_1499_3 ? _T_1548 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1550 = {auto_out_4_b_bits_id,auto_out_4_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1551 = _T_1499_4 ? _T_1550 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1552 = {auto_out_5_b_bits_id,auto_out_5_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1553 = _T_1499_5 ? _T_1552 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1554 = {auto_out_6_b_bits_id,auto_out_6_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1555 = _T_1499_6 ? _T_1554 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1556 = {auto_out_7_b_bits_id,auto_out_7_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1557 = _T_1499_7 ? _T_1556 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1558 = {auto_out_8_b_bits_id,auto_out_8_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1559 = _T_1499_8 ? _T_1558 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1560 = {auto_out_9_b_bits_id,auto_out_9_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1561 = _T_1499_9 ? _T_1560 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1562 = {auto_out_10_b_bits_id,auto_out_10_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1563 = _T_1499_10 ? _T_1562 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1564 = {auto_out_11_b_bits_id,auto_out_11_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1565 = _T_1499_11 ? _T_1564 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1566 = {auto_out_12_b_bits_id,auto_out_12_b_bits_resp}; // @[Mux.scala 27:72]
  assign _T_1567 = _T_1499_12 ? _T_1566 : 3'h0; // @[Mux.scala 27:72]
  assign _T_1568 = _T_1543 | _T_1545; // @[Mux.scala 27:72]
  assign _T_1569 = _T_1568 | _T_1547; // @[Mux.scala 27:72]
  assign _T_1570 = _T_1569 | _T_1549; // @[Mux.scala 27:72]
  assign _T_1571 = _T_1570 | _T_1551; // @[Mux.scala 27:72]
  assign _T_1572 = _T_1571 | _T_1553; // @[Mux.scala 27:72]
  assign _T_1573 = _T_1572 | _T_1555; // @[Mux.scala 27:72]
  assign _T_1574 = _T_1573 | _T_1557; // @[Mux.scala 27:72]
  assign _T_1575 = _T_1574 | _T_1559; // @[Mux.scala 27:72]
  assign _T_1576 = _T_1575 | _T_1561; // @[Mux.scala 27:72]
  assign _T_1577 = _T_1576 | _T_1563; // @[Mux.scala 27:72]
  assign _T_1578 = _T_1577 | _T_1565; // @[Mux.scala 27:72]
  assign _T_1579 = _T_1578 | _T_1567; // @[Mux.scala 27:72]
  assign auto_in_aw_ready = _T_268 & _T_260; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = in_0_w_ready & awIn_0_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = _T_1317 ? _T_1329 : _T_1539; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = _T_1579[1:0]; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = in_0_ar_ready & _T_232; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = _T_1022 ? _T_1034 : _T_1244; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = _T_1310[34:3]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = _T_1310[2:1]; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = _T_1310[0]; // @[LazyModule.scala 173:31]
  assign auto_out_12_aw_valid = in_0_aw_valid & requestAWIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_12_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_valid = in_0_w_valid & requestWIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_12_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_12_b_ready = auto_in_b_ready & _T_1501_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_valid = in_0_ar_valid & requestARIO_0_12; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_12_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_12_r_ready = auto_in_r_ready & _T_1206_12; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_valid = in_0_aw_valid & requestAWIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_11_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_valid = in_0_w_valid & requestWIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_11_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_11_b_ready = auto_in_b_ready & _T_1501_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_valid = in_0_ar_valid & requestARIO_0_11; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_11_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_11_r_ready = auto_in_r_ready & _T_1206_11; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_valid = in_0_aw_valid & requestAWIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_10_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_valid = in_0_w_valid & requestWIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_10_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_10_b_ready = auto_in_b_ready & _T_1501_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_valid = in_0_ar_valid & requestARIO_0_10; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_10_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_10_r_ready = auto_in_r_ready & _T_1206_10; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_valid = in_0_aw_valid & requestAWIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_9_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_valid = in_0_w_valid & requestWIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_9_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_9_b_ready = auto_in_b_ready & _T_1501_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_valid = in_0_ar_valid & requestARIO_0_9; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_9_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_9_r_ready = auto_in_r_ready & _T_1206_9; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_valid = in_0_aw_valid & requestAWIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_8_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_valid = in_0_w_valid & requestWIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_8_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_8_b_ready = auto_in_b_ready & _T_1501_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_valid = in_0_ar_valid & requestARIO_0_8; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_8_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_8_r_ready = auto_in_r_ready & _T_1206_8; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_valid = in_0_aw_valid & requestAWIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_7_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_valid = in_0_w_valid & requestWIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_7_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_7_b_ready = auto_in_b_ready & _T_1501_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_valid = in_0_ar_valid & requestARIO_0_7; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_7_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_7_r_ready = auto_in_r_ready & _T_1206_7; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_valid = in_0_aw_valid & requestAWIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_6_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_valid = in_0_w_valid & requestWIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_6_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_6_b_ready = auto_in_b_ready & _T_1501_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_valid = in_0_ar_valid & requestARIO_0_6; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_6_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_6_r_ready = auto_in_r_ready & _T_1206_6; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_valid = in_0_aw_valid & requestAWIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_5_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_valid = in_0_w_valid & requestWIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_5_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_5_b_ready = auto_in_b_ready & _T_1501_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_valid = in_0_ar_valid & requestARIO_0_5; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_5_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_5_r_ready = auto_in_r_ready & _T_1206_5; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_valid = in_0_aw_valid & requestAWIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_4_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_valid = in_0_w_valid & requestWIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_4_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_4_b_ready = auto_in_b_ready & _T_1501_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_valid = in_0_ar_valid & requestARIO_0_4; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_4_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_4_r_ready = auto_in_r_ready & _T_1206_4; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_valid = in_0_aw_valid & requestAWIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_3_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_valid = in_0_w_valid & requestWIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_3_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_3_b_ready = auto_in_b_ready & _T_1501_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_valid = in_0_ar_valid & requestARIO_0_3; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_3_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_3_r_ready = auto_in_r_ready & _T_1206_3; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_valid = in_0_aw_valid & requestAWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_valid = in_0_w_valid & requestWIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_2_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_2_b_ready = auto_in_b_ready & _T_1501_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_valid = in_0_ar_valid & requestARIO_0_2; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_2_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_2_r_ready = auto_in_r_ready & _T_1206_2; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_valid = in_0_aw_valid & requestAWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_valid = in_0_w_valid & requestWIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_1_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_1_b_ready = auto_in_b_ready & _T_1501_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_valid = in_0_ar_valid & requestARIO_0_1; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_1_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_1_r_ready = auto_in_r_ready & _T_1206_1; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_valid = in_0_aw_valid & requestAWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_addr = auto_in_aw_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_valid = in_0_w_valid & requestWIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_0_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_0_b_ready = auto_in_b_ready & _T_1501_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_valid = in_0_ar_valid & requestARIO_0_0; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_addr = auto_in_ar_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_0_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_0_r_ready = auto_in_r_ready & _T_1206_0; // @[LazyModule.scala 173:49]
  assign awIn_0_clock = clock;
  assign awIn_0_reset = reset;
  assign awIn_0_io_enq_valid = auto_in_aw_valid & _T_270; // @[Xbar.scala 140:30]
  assign awIn_0_io_enq_bits = {_T_140,_T_134}; // @[Xbar.scala 64:57]
  assign awIn_0_io_deq_ready = _T_276 & in_0_w_ready; // @[Xbar.scala 147:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_209 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_210 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1022 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1203_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1203_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1203_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1203_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1203_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1203_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1203_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1203_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1203_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1203_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1203_10 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1203_11 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1203_12 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1053 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_263 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_237 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_238 = _RAND_19[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1317 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1498_0 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1498_1 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1498_2 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1498_3 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1498_4 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1498_5 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1498_6 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1498_7 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1498_8 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_1498_9 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_1498_10 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1498_11 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_1498_12 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_1348 = _RAND_34[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_209 <= 3'h0;
    end else begin
      _T_209 <= _T_214;
    end
    if (_T_204) begin
      _T_210 <= _T_175;
    end
    _T_1022 <= reset | _GEN_58;
    if (reset) begin
      _T_1203_0 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_0 <= _T_1104;
    end
    if (reset) begin
      _T_1203_1 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_1 <= _T_1105;
    end
    if (reset) begin
      _T_1203_2 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_2 <= _T_1106;
    end
    if (reset) begin
      _T_1203_3 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_3 <= _T_1107;
    end
    if (reset) begin
      _T_1203_4 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_4 <= _T_1108;
    end
    if (reset) begin
      _T_1203_5 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_5 <= _T_1109;
    end
    if (reset) begin
      _T_1203_6 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_6 <= _T_1110;
    end
    if (reset) begin
      _T_1203_7 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_7 <= _T_1111;
    end
    if (reset) begin
      _T_1203_8 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_8 <= _T_1112;
    end
    if (reset) begin
      _T_1203_9 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_9 <= _T_1113;
    end
    if (reset) begin
      _T_1203_10 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_10 <= _T_1114;
    end
    if (reset) begin
      _T_1203_11 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_11 <= _T_1115;
    end
    if (reset) begin
      _T_1203_12 <= 1'h0;
    end else if (_T_1022) begin
      _T_1203_12 <= _T_1116;
    end
    if (reset) begin
      _T_1053 <= 13'h1fff;
    end else if (_T_1074) begin
      _T_1053 <= _T_1087;
    end
    if (reset) begin
      _T_263 <= 1'h0;
    end else if (_T_273) begin
      _T_263 <= 1'h0;
    end else begin
      _T_263 <= _GEN_2;
    end
    if (reset) begin
      _T_237 <= 3'h0;
    end else begin
      _T_237 <= _T_242;
    end
    if (_T_233) begin
      _T_238 <= _T_203;
    end
    _T_1317 <= reset | _GEN_61;
    if (reset) begin
      _T_1498_0 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_0 <= _T_1399;
    end
    if (reset) begin
      _T_1498_1 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_1 <= _T_1400;
    end
    if (reset) begin
      _T_1498_2 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_2 <= _T_1401;
    end
    if (reset) begin
      _T_1498_3 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_3 <= _T_1402;
    end
    if (reset) begin
      _T_1498_4 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_4 <= _T_1403;
    end
    if (reset) begin
      _T_1498_5 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_5 <= _T_1404;
    end
    if (reset) begin
      _T_1498_6 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_6 <= _T_1405;
    end
    if (reset) begin
      _T_1498_7 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_7 <= _T_1406;
    end
    if (reset) begin
      _T_1498_8 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_8 <= _T_1407;
    end
    if (reset) begin
      _T_1498_9 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_9 <= _T_1408;
    end
    if (reset) begin
      _T_1498_10 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_10 <= _T_1409;
    end
    if (reset) begin
      _T_1498_11 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_11 <= _T_1410;
    end
    if (reset) begin
      _T_1498_12 <= 1'h0;
    end else if (_T_1317) begin
      _T_1498_12 <= _T_1411;
    end
    if (reset) begin
      _T_1348 <= 13'h1fff;
    end else if (_T_1369) begin
      _T_1348 <= _T_1382;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_220) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_220) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_226) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_226) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_248) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:107 assert (!resp_fire || count =/= UInt(0))\n"); // @[Xbar.scala 107:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_248) begin
          $fatal; // @[Xbar.scala 107:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_254) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:108 assert (!req_fire  || count =/= UInt(flight))\n"); // @[Xbar.scala 108:22]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_254) begin
          $fatal; // @[Xbar.scala 108:22]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_465) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_465) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_486) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_486) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_509) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_509) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_530) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_530) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_553) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_553) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_574) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_574) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_597) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_597) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_618) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_618) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_641) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_641) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_662) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_662) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_685) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_685) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_706) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_706) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_729) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_729) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_750) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_750) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_773) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_773) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_794) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_794) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_817) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_817) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_838) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_838) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_861) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_861) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_882) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_882) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_905) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_905) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_926) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_926) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_949) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_949) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_970) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_970) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_993) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_993) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1014) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1014) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1184) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1184) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1201) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1479) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:256 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n"); // @[Xbar.scala 256:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1479) begin
          $fatal; // @[Xbar.scala 256:11]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1496) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Xbar.scala:258 assert (!anyValid || winner.reduce(_||_))\n"); // @[Xbar.scala 258:12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1496) begin
          $fatal; // @[Xbar.scala 258:12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_16(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [29:0] io_enq_bits_addr,
  input  [2:0]  io_enq_bits_size,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [29:0] io_deq_bits_addr,
  output [2:0]  io_deq_bits_size
);
  reg  _T_id [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 209:24]
  reg [29:0] _T_addr [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [29:0] _T_addr__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_18_addr; // @[Decoupled.scala 209:24]
  wire [29:0] _T_addr__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_addr__T_10_en; // @[Decoupled.scala 209:24]
  reg [2:0] _T_size [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [2:0] _T_size__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_size__T_18_addr; // @[Decoupled.scala 209:24]
  wire [2:0] _T_size__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_size__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_size__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_size__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_5;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_addr__T_18_addr = value_1;
  assign _T_addr__T_18_data = _T_addr[_T_addr__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_addr__T_10_data = io_enq_bits_addr;
  assign _T_addr__T_10_addr = value;
  assign _T_addr__T_10_mask = 1'h1;
  assign _T_addr__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_size__T_18_addr = value_1;
  assign _T_size__T_18_data = _T_size[_T_size__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_size__T_10_data = io_enq_bits_size;
  assign _T_size__T_10_addr = value;
  assign _T_size__T_10_mask = 1'h1;
  assign _T_size__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_addr = _T_addr__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_size = _T_size__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_addr[initvar] = _RAND_1[29:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_addr__T_10_en & _T_addr__T_10_mask) begin
      _T_addr[_T_addr__T_10_addr] <= _T_addr__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_size__T_10_en & _T_size__T_10_mask) begin
      _T_size[_T_size__T_10_addr] <= _T_size__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input  [3:0]  io_enq_bits_strb,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output [3:0]  io_deq_bits_strb
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg [3:0] _T_strb [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [3:0] _T_strb__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_18_addr; // @[Decoupled.scala 209:24]
  wire [3:0] _T_strb__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_strb__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_strb__T_18_addr = value_1;
  assign _T_strb__T_18_data = _T_strb[_T_strb__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_strb__T_10_data = io_enq_bits_strb;
  assign _T_strb__T_10_addr = value;
  assign _T_strb__T_10_mask = 1'h1;
  assign _T_strb__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_strb = _T_strb__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_strb[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_strb__T_10_en & _T_strb__T_10_mask) begin
      _T_strb[_T_strb__T_10_addr] <= _T_strb__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_18(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg  _T_id [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] _T_resp [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [1:0] _T_resp__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_18_addr; // @[Decoupled.scala 209:24]
  wire [1:0] _T_resp__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_resp__T_10_data = 2'h0;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_resp = _T_resp__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module Queue_20(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg  _T_id [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire  _T_id__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 209:24]
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg [1:0] _T_resp [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_2;
  wire [1:0] _T_resp__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_18_addr; // @[Decoupled.scala 209:24]
  wire [1:0] _T_resp__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_resp__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_3;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_6;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_id__T_18_addr = value_1;
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_resp__T_18_addr = value_1;
  assign _T_resp__T_18_data = _T_resp[_T_resp__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_resp__T_10_data = 2'h0;
  assign _T_resp__T_10_addr = value;
  assign _T_resp__T_10_mask = 1'h1;
  assign _T_resp__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = 1'h1;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_resp = _T_resp__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_resp__T_10_en & _T_resp__T_10_mask) begin
      _T_resp[_T_resp__T_10_addr] <= _T_resp__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4Buffer(
  input         clock,
  input         reset,
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [29:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output        auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [29:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output        auto_in_r_bits_id,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input         auto_out_b_bits_id,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input         auto_out_r_bits_id,
  input  [31:0] auto_out_r_bits_data
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_io_enq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_io_enq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_io_deq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_io_deq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_1_clock; // @[Decoupled.scala 287:21]
  wire  Queue_1_reset; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_1_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire [3:0] Queue_1_io_enq_bits_strb; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_1_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_1_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire [3:0] Queue_1_io_deq_bits_strb; // @[Decoupled.scala 287:21]
  wire  Queue_2_clock; // @[Decoupled.scala 287:21]
  wire  Queue_2_reset; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_2_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [1:0] Queue_2_io_deq_bits_resp; // @[Decoupled.scala 287:21]
  wire  Queue_3_clock; // @[Decoupled.scala 287:21]
  wire  Queue_3_reset; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_3_io_enq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_3_io_enq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_3_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [29:0] Queue_3_io_deq_bits_addr; // @[Decoupled.scala 287:21]
  wire [2:0] Queue_3_io_deq_bits_size; // @[Decoupled.scala 287:21]
  wire  Queue_4_clock; // @[Decoupled.scala 287:21]
  wire  Queue_4_reset; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_enq_bits_id; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_4_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_valid; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_bits_id; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_4_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire [1:0] Queue_4_io_deq_bits_resp; // @[Decoupled.scala 287:21]
  wire  Queue_4_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_16 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_size(Queue_io_deq_bits_size)
  );
  Queue_17 Queue_1 ( // @[Decoupled.scala 287:21]
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb)
  );
  Queue_18 Queue_2 ( // @[Decoupled.scala 287:21]
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  Queue_16 Queue_3 ( // @[Decoupled.scala 287:21]
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_size(Queue_3_io_deq_bits_size)
  );
  Queue_20 Queue_4 ( // @[Decoupled.scala 287:21]
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign auto_in_aw_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = Queue_1_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = Queue_2_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_id = Queue_2_io_deq_bits_id; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = Queue_2_io_deq_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = Queue_3_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = Queue_4_io_deq_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_id = Queue_4_io_deq_bits_id; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = Queue_4_io_deq_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = Queue_4_io_deq_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = Queue_4_io_deq_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = Queue_io_deq_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = Queue_io_deq_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = Queue_1_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = Queue_1_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = Queue_1_io_deq_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = Queue_2_io_enq_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = Queue_3_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = Queue_3_io_deq_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = Queue_3_io_deq_bits_addr; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = Queue_3_io_deq_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = Queue_4_io_enq_ready; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_aw_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_id = auto_in_aw_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_addr = auto_in_aw_bits_addr; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_size = auto_in_aw_bits_size; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_aw_ready; // @[Decoupled.scala 311:15]
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = auto_in_w_valid; // @[Decoupled.scala 288:22]
  assign Queue_1_io_enq_bits_data = auto_in_w_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_1_io_enq_bits_strb = auto_in_w_bits_strb; // @[Decoupled.scala 289:21]
  assign Queue_1_io_deq_ready = auto_out_w_ready; // @[Decoupled.scala 311:15]
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = auto_out_b_valid; // @[Decoupled.scala 288:22]
  assign Queue_2_io_enq_bits_id = auto_out_b_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_2_io_deq_ready = auto_in_b_ready; // @[Decoupled.scala 311:15]
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = auto_in_ar_valid; // @[Decoupled.scala 288:22]
  assign Queue_3_io_enq_bits_id = auto_in_ar_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_3_io_enq_bits_addr = auto_in_ar_bits_addr; // @[Decoupled.scala 289:21]
  assign Queue_3_io_enq_bits_size = auto_in_ar_bits_size; // @[Decoupled.scala 289:21]
  assign Queue_3_io_deq_ready = auto_out_ar_ready; // @[Decoupled.scala 311:15]
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = auto_out_r_valid; // @[Decoupled.scala 288:22]
  assign Queue_4_io_enq_bits_id = auto_out_r_bits_id; // @[Decoupled.scala 289:21]
  assign Queue_4_io_enq_bits_data = auto_out_r_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_4_io_deq_ready = auto_in_r_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_81(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_81 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_88(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_7(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_88 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module Queue_97(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_last
);
  reg [31:0] _T_data [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_0;
  wire [31:0] _T_data__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_18_addr; // @[Decoupled.scala 209:24]
  wire [31:0] _T_data__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_data__T_10_en; // @[Decoupled.scala 209:24]
  reg  _T_last [0:1]; // @[Decoupled.scala 209:24]
  reg [31:0] _RAND_1;
  wire  _T_last__T_18_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_18_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_data; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_addr; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_mask; // @[Decoupled.scala 209:24]
  wire  _T_last__T_10_en; // @[Decoupled.scala 209:24]
  reg  value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_2;
  reg  value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  reg  _T_1; // @[Decoupled.scala 212:35]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 214:41]
  wire  _T_3; // @[Decoupled.scala 215:36]
  wire  _T_4; // @[Decoupled.scala 215:33]
  wire  _T_5; // @[Decoupled.scala 216:32]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Counter.scala 39:22]
  wire  _T_14; // @[Counter.scala 39:22]
  wire  _T_15; // @[Decoupled.scala 227:16]
  assign _T_data__T_18_addr = value_1;
  assign _T_data__T_18_data = _T_data[_T_data__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_data__T_10_data = io_enq_bits_data;
  assign _T_data__T_10_addr = value;
  assign _T_data__T_10_mask = 1'h1;
  assign _T_data__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_last__T_18_addr = value_1;
  assign _T_last__T_18_data = _T_last[_T_last__T_18_addr]; // @[Decoupled.scala 209:24]
  assign _T_last__T_10_data = io_enq_bits_last;
  assign _T_last__T_10_addr = value;
  assign _T_last__T_10_mask = 1'h1;
  assign _T_last__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_2 = value == value_1; // @[Decoupled.scala 214:41]
  assign _T_3 = ~_T_1; // @[Decoupled.scala 215:36]
  assign _T_4 = _T_2 & _T_3; // @[Decoupled.scala 215:33]
  assign _T_5 = _T_2 & _T_1; // @[Decoupled.scala 216:32]
  assign _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = value + 1'h1; // @[Counter.scala 39:22]
  assign _T_14 = value_1 + 1'h1; // @[Counter.scala 39:22]
  assign _T_15 = _T_6 != _T_8; // @[Decoupled.scala 227:16]
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 232:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 231:16]
  assign io_deq_bits_data = _T_data__T_18_data; // @[Decoupled.scala 233:15]
  assign io_deq_bits_last = _T_last__T_18_data; // @[Decoupled.scala 233:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_data[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    _T_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_data__T_10_en & _T_data__T_10_mask) begin
      _T_data[_T_data__T_10_addr] <= _T_data__T_10_data; // @[Decoupled.scala 209:24]
    end
    if(_T_last__T_10_en & _T_last__T_10_mask) begin
      _T_last[_T_last__T_10_addr] <= _T_last__T_10_data; // @[Decoupled.scala 209:24]
    end
    if (reset) begin
      value <= 1'h0;
    end else if (_T_6) begin
      value <= _T_12;
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else if (_T_8) begin
      value_1 <= _T_14;
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module AXI4StreamBuffer_16(
  input         clock,
  input         reset,
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  wire  Queue_clock; // @[Decoupled.scala 287:21]
  wire  Queue_reset; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_enq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_enq_bits_last; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_ready; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_valid; // @[Decoupled.scala 287:21]
  wire [31:0] Queue_io_deq_bits_data; // @[Decoupled.scala 287:21]
  wire  Queue_io_deq_bits_last; // @[Decoupled.scala 287:21]
  Queue_97 Queue ( // @[Decoupled.scala 287:21]
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  assign auto_in_ready = Queue_io_enq_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = Queue_io_deq_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = Queue_io_deq_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = Queue_io_deq_bits_last; // @[LazyModule.scala 173:49]
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = auto_in_valid; // @[Decoupled.scala 288:22]
  assign Queue_io_enq_bits_data = auto_in_bits_data; // @[Decoupled.scala 289:21]
  assign Queue_io_enq_bits_last = auto_in_bits_last; // @[Decoupled.scala 289:21]
  assign Queue_io_deq_ready = auto_out_ready; // @[Decoupled.scala 311:15]
endmodule
module BundleBridgeToAXI4(
  output        auto_in_aw_ready,
  input         auto_in_aw_valid,
  input         auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [2:0]  auto_in_aw_bits_size,
  output        auto_in_w_ready,
  input         auto_in_w_valid,
  input  [31:0] auto_in_w_bits_data,
  input  [3:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
  input         auto_in_b_ready,
  output        auto_in_b_valid,
  output [1:0]  auto_in_b_bits_resp,
  output        auto_in_ar_ready,
  input         auto_in_ar_valid,
  input         auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [2:0]  auto_in_ar_bits_size,
  input         auto_in_r_ready,
  output        auto_in_r_valid,
  output [31:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output        auto_in_r_bits_last,
  input         auto_out_aw_ready,
  output        auto_out_aw_valid,
  output        auto_out_aw_bits_id,
  output [29:0] auto_out_aw_bits_addr,
  output [2:0]  auto_out_aw_bits_size,
  input         auto_out_w_ready,
  output        auto_out_w_valid,
  output [31:0] auto_out_w_bits_data,
  output [3:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
  output        auto_out_b_ready,
  input         auto_out_b_valid,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
  output        auto_out_ar_valid,
  output        auto_out_ar_bits_id,
  output [29:0] auto_out_ar_bits_addr,
  output [2:0]  auto_out_ar_bits_size,
  output        auto_out_r_ready,
  input         auto_out_r_valid,
  input  [31:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last
);
  assign auto_in_aw_ready = auto_out_aw_ready; // @[LazyModule.scala 173:31]
  assign auto_in_w_ready = auto_out_w_ready; // @[LazyModule.scala 173:31]
  assign auto_in_b_valid = auto_out_b_valid; // @[LazyModule.scala 173:31]
  assign auto_in_b_bits_resp = auto_out_b_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_ar_ready = auto_out_ar_ready; // @[LazyModule.scala 173:31]
  assign auto_in_r_valid = auto_out_r_valid; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_data = auto_out_r_bits_data; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_resp = auto_out_r_bits_resp; // @[LazyModule.scala 173:31]
  assign auto_in_r_bits_last = auto_out_r_bits_last; // @[LazyModule.scala 173:31]
  assign auto_out_aw_valid = auto_in_aw_valid; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_id = auto_in_aw_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_aw_bits_size = auto_in_aw_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_w_valid = auto_in_w_valid; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_data = auto_in_w_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_strb = auto_in_w_bits_strb; // @[LazyModule.scala 173:49]
  assign auto_out_w_bits_last = auto_in_w_bits_last; // @[LazyModule.scala 173:49]
  assign auto_out_b_ready = auto_in_b_ready; // @[LazyModule.scala 173:49]
  assign auto_out_ar_valid = auto_in_ar_valid; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_id = auto_in_ar_bits_id; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr[29:0]; // @[LazyModule.scala 173:49]
  assign auto_out_ar_bits_size = auto_in_ar_bits_size; // @[LazyModule.scala 173:49]
  assign auto_out_r_ready = auto_in_r_ready; // @[LazyModule.scala 173:49]
endmodule
module AXI4StreamToBundleBridge(
  output       auto_in_ready,
  input        auto_in_valid,
  input  [7:0] auto_in_bits_data,
  input        auto_in_bits_last,
  input        auto_out_ready,
  output       auto_out_valid,
  output [7:0] auto_out_bits_data,
  output       auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module AXI4StreamToBundleBridge_1(
  output        auto_in_ready,
  input         auto_in_valid,
  input  [31:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [31:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module LISTestWithLA(
  input         clock,
  input         reset,
  output        ioMem_0_aw_ready,
  input         ioMem_0_aw_valid,
  input         ioMem_0_aw_bits_id,
  input  [31:0] ioMem_0_aw_bits_addr,
  input  [7:0]  ioMem_0_aw_bits_len,
  input  [2:0]  ioMem_0_aw_bits_size,
  input  [1:0]  ioMem_0_aw_bits_burst,
  input         ioMem_0_aw_bits_lock,
  input  [3:0]  ioMem_0_aw_bits_cache,
  input  [2:0]  ioMem_0_aw_bits_prot,
  input  [3:0]  ioMem_0_aw_bits_qos,
  output        ioMem_0_w_ready,
  input         ioMem_0_w_valid,
  input  [31:0] ioMem_0_w_bits_data,
  input  [3:0]  ioMem_0_w_bits_strb,
  input         ioMem_0_w_bits_last,
  input         ioMem_0_b_ready,
  output        ioMem_0_b_valid,
  output        ioMem_0_b_bits_id,
  output [1:0]  ioMem_0_b_bits_resp,
  output        ioMem_0_ar_ready,
  input         ioMem_0_ar_valid,
  input         ioMem_0_ar_bits_id,
  input  [31:0] ioMem_0_ar_bits_addr,
  input  [7:0]  ioMem_0_ar_bits_len,
  input  [2:0]  ioMem_0_ar_bits_size,
  input  [1:0]  ioMem_0_ar_bits_burst,
  input         ioMem_0_ar_bits_lock,
  input  [3:0]  ioMem_0_ar_bits_cache,
  input  [2:0]  ioMem_0_ar_bits_prot,
  input  [3:0]  ioMem_0_ar_bits_qos,
  input         ioMem_0_r_ready,
  output        ioMem_0_r_valid,
  output        ioMem_0_r_bits_id,
  output [31:0] ioMem_0_r_bits_data,
  output [1:0]  ioMem_0_r_bits_resp,
  output        ioMem_0_r_bits_last,
  input         outStream_0_ready,
  output        outStream_0_valid,
  output [7:0]  outStream_0_bits_data,
  output        outStream_0_bits_last,
  output        inStream_0_ready,
  input         inStream_0_valid,
  input  [7:0]  inStream_0_bits_data,
  input         inStream_0_bits_last,
  input         laInside_0_ready,
  output        laInside_0_valid,
  output [31:0] laInside_0_bits_data,
  output        laInside_0_bits_last,
  input         laOutside_0_ready,
  output        laOutside_0_valid,
  output [31:0] laOutside_0_bits_data,
  output        laOutside_0_bits_last,
  output        int_0,
  output        uTx,
  input         uRx
);
  wire  widthAdapter_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  in_split_clock; // @[LISTestWithLA.scala 55:29]
  wire  in_split_reset; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 55:29]
  wire [29:0] in_split_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_w_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_w_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 55:29]
  wire [3:0] in_split_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_b_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_b_valid; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 55:29]
  wire [29:0] in_split_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 55:29]
  wire [2:0] in_split_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_r_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_r_valid; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_in_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_in_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_stream_in_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_in_bits_last; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_4_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_4_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_stream_out_4_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_4_bits_last; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_3_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_3_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_stream_out_3_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_3_bits_last; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_2_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_2_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_stream_out_2_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_2_bits_last; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_1_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_1_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_stream_out_1_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_1_bits_last; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_0_ready; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_0_valid; // @[LISTestWithLA.scala 55:29]
  wire [31:0] in_split_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 55:29]
  wire  in_split_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 55:29]
  wire  in_queue_clock; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_reset; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_auto_out_out_ready; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_auto_out_out_valid; // @[LISTestWithLA.scala 56:29]
  wire [7:0] in_queue_auto_out_out_bits_data; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_auto_out_out_bits_last; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_auto_in_in_ready; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_auto_in_in_valid; // @[LISTestWithLA.scala 56:29]
  wire [7:0] in_queue_auto_in_in_bits_data; // @[LISTestWithLA.scala 56:29]
  wire  in_queue_auto_in_in_bits_last; // @[LISTestWithLA.scala 56:29]
  wire  lisFifo_clock; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_reset; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 59:33]
  wire [29:0] lisFifo_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_w_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_w_valid; // @[LISTestWithLA.scala 59:33]
  wire [31:0] lisFifo_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 59:33]
  wire [3:0] lisFifo_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_b_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_b_valid; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 59:33]
  wire [29:0] lisFifo_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 59:33]
  wire [2:0] lisFifo_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_r_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_r_valid; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 59:33]
  wire [31:0] lisFifo_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_stream_in_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_stream_in_valid; // @[LISTestWithLA.scala 59:33]
  wire [31:0] lisFifo_auto_stream_in_bits_data; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_stream_in_bits_last; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_stream_out_ready; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_stream_out_valid; // @[LISTestWithLA.scala 59:33]
  wire [31:0] lisFifo_auto_stream_out_bits_data; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_auto_stream_out_bits_last; // @[LISTestWithLA.scala 59:33]
  wire  lisFifo_mux0_clock; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_reset; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_aw_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_aw_valid; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_aw_bits_id; // @[LISTestWithLA.scala 60:33]
  wire [29:0] lisFifo_mux0_auto_register_in_aw_bits_addr; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_w_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_w_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_register_in_w_bits_data; // @[LISTestWithLA.scala 60:33]
  wire [3:0] lisFifo_mux0_auto_register_in_w_bits_strb; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_b_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_b_valid; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_b_bits_id; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_ar_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_ar_valid; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_ar_bits_id; // @[LISTestWithLA.scala 60:33]
  wire [29:0] lisFifo_mux0_auto_register_in_ar_bits_addr; // @[LISTestWithLA.scala 60:33]
  wire [2:0] lisFifo_mux0_auto_register_in_ar_bits_size; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_r_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_r_valid; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_register_in_r_bits_id; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_register_in_r_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_4_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_4_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_stream_in_4_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_4_bits_last; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_3_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_3_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_stream_in_3_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_3_bits_last; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_2_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_2_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_stream_in_2_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_2_bits_last; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_1_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_1_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_stream_in_1_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_1_bits_last; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_0_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_0_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_stream_in_0_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_in_0_bits_last; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_out_0_ready; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_out_0_valid; // @[LISTestWithLA.scala 60:33]
  wire [31:0] lisFifo_mux0_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 60:33]
  wire  lisFifo_mux0_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 60:33]
  wire  lisInput_clock; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_reset; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 66:34]
  wire [29:0] lisInput_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_w_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_w_valid; // @[LISTestWithLA.scala 66:34]
  wire [31:0] lisInput_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 66:34]
  wire [3:0] lisInput_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_b_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_b_valid; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 66:34]
  wire [29:0] lisInput_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 66:34]
  wire [2:0] lisInput_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_r_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_r_valid; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 66:34]
  wire [31:0] lisInput_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_stream_in_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_stream_in_valid; // @[LISTestWithLA.scala 66:34]
  wire [31:0] lisInput_auto_stream_in_bits_data; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_stream_in_bits_last; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_stream_out_ready; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_stream_out_valid; // @[LISTestWithLA.scala 66:34]
  wire [31:0] lisInput_auto_stream_out_bits_data; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_auto_stream_out_bits_last; // @[LISTestWithLA.scala 66:34]
  wire  lisInput_mux0_clock; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_reset; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_aw_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_aw_valid; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_aw_bits_id; // @[LISTestWithLA.scala 67:34]
  wire [29:0] lisInput_mux0_auto_register_in_aw_bits_addr; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_w_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_w_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_register_in_w_bits_data; // @[LISTestWithLA.scala 67:34]
  wire [3:0] lisInput_mux0_auto_register_in_w_bits_strb; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_b_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_b_valid; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_b_bits_id; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_ar_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_ar_valid; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_ar_bits_id; // @[LISTestWithLA.scala 67:34]
  wire [29:0] lisInput_mux0_auto_register_in_ar_bits_addr; // @[LISTestWithLA.scala 67:34]
  wire [2:0] lisInput_mux0_auto_register_in_ar_bits_size; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_r_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_r_valid; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_register_in_r_bits_id; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_register_in_r_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_4_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_4_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_stream_in_4_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_4_bits_last; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_3_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_3_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_stream_in_3_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_3_bits_last; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_2_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_2_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_stream_in_2_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_2_bits_last; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_1_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_1_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_stream_in_1_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_1_bits_last; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_0_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_0_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_stream_in_0_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_in_0_bits_last; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_out_0_ready; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_out_0_valid; // @[LISTestWithLA.scala 67:34]
  wire [31:0] lisInput_mux0_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 67:34]
  wire  lisInput_mux0_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 67:34]
  wire  lisFixed_clock; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_reset; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 73:34]
  wire [29:0] lisFixed_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_w_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_w_valid; // @[LISTestWithLA.scala 73:34]
  wire [31:0] lisFixed_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 73:34]
  wire [3:0] lisFixed_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_b_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_b_valid; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 73:34]
  wire [29:0] lisFixed_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 73:34]
  wire [2:0] lisFixed_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_r_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_r_valid; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 73:34]
  wire [31:0] lisFixed_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_stream_in_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_stream_in_valid; // @[LISTestWithLA.scala 73:34]
  wire [31:0] lisFixed_auto_stream_in_bits_data; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_stream_in_bits_last; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_stream_out_ready; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_stream_out_valid; // @[LISTestWithLA.scala 73:34]
  wire [31:0] lisFixed_auto_stream_out_bits_data; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_auto_stream_out_bits_last; // @[LISTestWithLA.scala 73:34]
  wire  lisFixed_mux0_clock; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_reset; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_aw_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_aw_valid; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_aw_bits_id; // @[LISTestWithLA.scala 74:34]
  wire [29:0] lisFixed_mux0_auto_register_in_aw_bits_addr; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_w_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_w_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_register_in_w_bits_data; // @[LISTestWithLA.scala 74:34]
  wire [3:0] lisFixed_mux0_auto_register_in_w_bits_strb; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_b_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_b_valid; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_b_bits_id; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_ar_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_ar_valid; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_ar_bits_id; // @[LISTestWithLA.scala 74:34]
  wire [29:0] lisFixed_mux0_auto_register_in_ar_bits_addr; // @[LISTestWithLA.scala 74:34]
  wire [2:0] lisFixed_mux0_auto_register_in_ar_bits_size; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_r_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_r_valid; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_register_in_r_bits_id; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_register_in_r_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_4_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_4_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_stream_in_4_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_4_bits_last; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_3_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_3_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_stream_in_3_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_3_bits_last; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_2_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_2_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_stream_in_2_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_2_bits_last; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_1_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_1_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_stream_in_1_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_1_bits_last; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_0_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_0_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_stream_in_0_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_in_0_bits_last; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_out_0_ready; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_out_0_valid; // @[LISTestWithLA.scala 74:34]
  wire [31:0] lisFixed_mux0_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 74:34]
  wire  lisFixed_mux0_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 74:34]
  wire  bist_clock; // @[LISTestWithLA.scala 79:34]
  wire  bist_reset; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 79:34]
  wire [29:0] bist_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_w_ready; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_w_valid; // @[LISTestWithLA.scala 79:34]
  wire [31:0] bist_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 79:34]
  wire [3:0] bist_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_b_ready; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_b_valid; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 79:34]
  wire [29:0] bist_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 79:34]
  wire [2:0] bist_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_r_ready; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_r_valid; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 79:34]
  wire [31:0] bist_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_stream_out_ready; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_stream_out_valid; // @[LISTestWithLA.scala 79:34]
  wire [31:0] bist_auto_stream_out_bits_data; // @[LISTestWithLA.scala 79:34]
  wire  bist_auto_stream_out_bits_last; // @[LISTestWithLA.scala 79:34]
  wire  bist_split_clock; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_reset; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 80:34]
  wire [29:0] bist_split_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_w_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_w_valid; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 80:34]
  wire [3:0] bist_split_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_b_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_b_valid; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 80:34]
  wire [29:0] bist_split_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 80:34]
  wire [2:0] bist_split_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_r_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_r_valid; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_in_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_in_valid; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_stream_in_bits_data; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_in_bits_last; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_3_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_3_valid; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_stream_out_3_bits_data; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_3_bits_last; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_2_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_2_valid; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_stream_out_2_bits_data; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_2_bits_last; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_1_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_1_valid; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_stream_out_1_bits_data; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_1_bits_last; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_0_ready; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_0_valid; // @[LISTestWithLA.scala 80:34]
  wire [31:0] bist_split_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 80:34]
  wire  bist_split_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 80:34]
  wire  out_mux_clock; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_reset; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_aw_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_aw_valid; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_aw_bits_id; // @[LISTestWithLA.scala 83:29]
  wire [29:0] out_mux_auto_register_in_aw_bits_addr; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_w_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_w_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_register_in_w_bits_data; // @[LISTestWithLA.scala 83:29]
  wire [3:0] out_mux_auto_register_in_w_bits_strb; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_b_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_b_valid; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_b_bits_id; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_ar_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_ar_valid; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_ar_bits_id; // @[LISTestWithLA.scala 83:29]
  wire [29:0] out_mux_auto_register_in_ar_bits_addr; // @[LISTestWithLA.scala 83:29]
  wire [2:0] out_mux_auto_register_in_ar_bits_size; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_r_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_r_valid; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_register_in_r_bits_id; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_register_in_r_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_5_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_5_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_in_5_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_5_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_4_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_4_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_in_4_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_4_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_3_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_3_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_in_3_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_3_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_2_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_2_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_in_2_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_2_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_1_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_1_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_in_1_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_1_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_0_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_0_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_in_0_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_in_0_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_out_1_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_out_1_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_out_1_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_out_1_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_out_0_ready; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_out_0_valid; // @[LISTestWithLA.scala 83:29]
  wire [31:0] out_mux_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 83:29]
  wire  out_mux_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 83:29]
  wire  out_split_clock; // @[LISTestWithLA.scala 84:29]
  wire  out_split_reset; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 84:29]
  wire [29:0] out_split_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_w_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_w_valid; // @[LISTestWithLA.scala 84:29]
  wire [31:0] out_split_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 84:29]
  wire [3:0] out_split_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_b_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_b_valid; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 84:29]
  wire [29:0] out_split_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 84:29]
  wire [2:0] out_split_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_r_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_r_valid; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 84:29]
  wire [31:0] out_split_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_in_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_in_valid; // @[LISTestWithLA.scala 84:29]
  wire [31:0] out_split_auto_stream_in_bits_data; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_in_bits_last; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_out_1_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_out_1_valid; // @[LISTestWithLA.scala 84:29]
  wire [31:0] out_split_auto_stream_out_1_bits_data; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_out_1_bits_last; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_out_0_ready; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_out_0_valid; // @[LISTestWithLA.scala 84:29]
  wire [31:0] out_split_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 84:29]
  wire  out_split_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 84:29]
  wire  out_queue_clock; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_reset; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_auto_out_out_ready; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_auto_out_out_valid; // @[LISTestWithLA.scala 85:29]
  wire [31:0] out_queue_auto_out_out_bits_data; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_auto_out_out_bits_last; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_auto_in_in_ready; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_auto_in_in_valid; // @[LISTestWithLA.scala 85:29]
  wire [31:0] out_queue_auto_in_in_bits_data; // @[LISTestWithLA.scala 85:29]
  wire  out_queue_auto_in_in_bits_last; // @[LISTestWithLA.scala 85:29]
  wire  widthAdapter_1_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_1_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_1_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_1_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  uTx_queue_clock; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_reset; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_auto_out_out_ready; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_auto_out_out_valid; // @[LISTestWithLA.scala 89:29]
  wire [31:0] uTx_queue_auto_out_out_bits_data; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_auto_out_out_bits_last; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_auto_in_in_ready; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_auto_in_in_valid; // @[LISTestWithLA.scala 89:29]
  wire [31:0] uTx_queue_auto_in_in_bits_data; // @[LISTestWithLA.scala 89:29]
  wire  uTx_queue_auto_in_in_bits_last; // @[LISTestWithLA.scala 89:29]
  wire  widthAdapter_2_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_2_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_in_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_2_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_2_auto_out_bits_last; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_clock; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_reset; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_in_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [7:0] widthAdapter_3_auto_in_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_ready; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  widthAdapter_3_auto_out_valid; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire [31:0] widthAdapter_3_auto_out_bits_data; // @[AXI4StreamWidthAdapter.scala 82:34]
  wire  uRx_split_clock; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_reset; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 92:29]
  wire [29:0] uRx_split_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_w_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_w_valid; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 92:29]
  wire [3:0] uRx_split_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_b_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_b_valid; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 92:29]
  wire [29:0] uRx_split_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 92:29]
  wire [2:0] uRx_split_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_r_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_r_valid; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_in_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_in_valid; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_stream_in_bits_data; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_in_bits_last; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_3_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_3_valid; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_stream_out_3_bits_data; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_3_bits_last; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_2_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_2_valid; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_stream_out_2_bits_data; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_2_bits_last; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_1_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_1_valid; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_stream_out_1_bits_data; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_1_bits_last; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_0_ready; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_0_valid; // @[LISTestWithLA.scala 92:29]
  wire [31:0] uRx_split_auto_stream_out_0_bits_data; // @[LISTestWithLA.scala 92:29]
  wire  uRx_split_auto_stream_out_0_bits_last; // @[LISTestWithLA.scala 92:29]
  wire  uart_clock; // @[LISTestWithLA.scala 93:29]
  wire  uart_reset; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_aw_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_aw_valid; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_aw_bits_id; // @[LISTestWithLA.scala 93:29]
  wire [29:0] uart_auto_mem_in_aw_bits_addr; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_w_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_w_valid; // @[LISTestWithLA.scala 93:29]
  wire [31:0] uart_auto_mem_in_w_bits_data; // @[LISTestWithLA.scala 93:29]
  wire [3:0] uart_auto_mem_in_w_bits_strb; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_b_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_b_valid; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_b_bits_id; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_ar_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_ar_valid; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_ar_bits_id; // @[LISTestWithLA.scala 93:29]
  wire [29:0] uart_auto_mem_in_ar_bits_addr; // @[LISTestWithLA.scala 93:29]
  wire [2:0] uart_auto_mem_in_ar_bits_size; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_r_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_r_valid; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_mem_in_r_bits_id; // @[LISTestWithLA.scala 93:29]
  wire [31:0] uart_auto_mem_in_r_bits_data; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_in_in_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_in_in_valid; // @[LISTestWithLA.scala 93:29]
  wire [7:0] uart_auto_in_in_bits_data; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_out_out_ready; // @[LISTestWithLA.scala 93:29]
  wire  uart_auto_out_out_valid; // @[LISTestWithLA.scala 93:29]
  wire [7:0] uart_auto_out_out_bits_data; // @[LISTestWithLA.scala 93:29]
  wire  uart_int_0; // @[LISTestWithLA.scala 93:29]
  wire  uart_io_txd; // @[LISTestWithLA.scala 93:29]
  wire  uart_io_rxd; // @[LISTestWithLA.scala 93:29]
  wire  bus_clock; // @[LISTestWithLA.scala 108:23]
  wire  bus_reset; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_in_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_in_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_in_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_in_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_w_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_b_valid; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_in_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_in_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_in_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_r_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_in_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_in_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_in_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_12_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_12_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_12_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_12_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_12_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_12_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_12_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_12_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_12_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_12_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_11_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_11_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_11_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_11_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_11_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_11_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_11_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_11_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_11_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_11_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_10_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_10_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_10_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_10_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_10_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_10_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_10_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_10_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_10_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_10_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_9_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_9_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_9_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_9_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_9_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_9_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_9_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_9_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_9_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_9_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_8_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_8_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_8_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_8_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_8_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_8_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_8_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_8_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_8_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_8_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_7_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_7_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_7_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_7_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_7_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_7_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_7_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_7_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_7_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_7_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_6_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_6_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_6_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_6_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_6_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_6_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_6_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_6_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_6_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_6_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_5_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_5_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_5_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_5_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_5_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_5_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_5_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_5_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_5_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_5_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_4_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_4_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_4_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_4_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_4_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_4_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_4_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_4_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_4_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_4_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_3_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_3_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_3_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_3_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_3_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_3_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_3_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_3_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_3_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_3_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_2_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_2_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_2_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_2_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_2_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_2_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_2_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_2_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_2_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_2_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_1_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_1_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_1_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_1_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_1_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_1_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_1_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_1_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_1_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_1_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_aw_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_aw_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_aw_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_0_aw_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_0_aw_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_w_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_w_valid; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_0_w_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [3:0] bus_auto_out_0_w_bits_strb; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_b_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_b_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_b_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_0_b_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_ar_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_ar_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_ar_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [29:0] bus_auto_out_0_ar_bits_addr; // @[LISTestWithLA.scala 108:23]
  wire [2:0] bus_auto_out_0_ar_bits_size; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_r_ready; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_r_valid; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_r_bits_id; // @[LISTestWithLA.scala 108:23]
  wire [31:0] bus_auto_out_0_r_bits_data; // @[LISTestWithLA.scala 108:23]
  wire [1:0] bus_auto_out_0_r_bits_resp; // @[LISTestWithLA.scala 108:23]
  wire  bus_auto_out_0_r_bits_last; // @[LISTestWithLA.scala 108:23]
  wire  axi4buf_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_1_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_1_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_1_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_1_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_1_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_1_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_1_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_1_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_2_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_2_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_2_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_2_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_2_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_2_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_2_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_2_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_2_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_3_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_3_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_3_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_3_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_3_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_3_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_3_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_3_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_3_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_4_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_4_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_4_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_4_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_4_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_4_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_4_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_4_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_4_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_5_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_5_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_5_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_5_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_5_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_5_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_5_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_5_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_5_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_6_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_6_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_6_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_6_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_6_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_6_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_6_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_6_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_6_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_7_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_7_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_7_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_7_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_7_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_7_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_7_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_7_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_7_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_8_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_8_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_8_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_8_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_8_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_8_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_8_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_8_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_8_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_9_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_9_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_9_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_9_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_9_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_9_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_9_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_9_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_9_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_10_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_10_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_10_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_10_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_10_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_10_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_10_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_10_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_10_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_11_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_11_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_11_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_11_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_11_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_11_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_11_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_11_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_11_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  axi4buf_12_clock; // @[Buffer.scala 58:29]
  wire  axi4buf_12_reset; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_in_aw_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_in_aw_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_in_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_12_auto_in_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_b_bits_id; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_in_b_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_in_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_in_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_in_r_bits_data; // @[Buffer.scala 58:29]
  wire [1:0] axi4buf_12_auto_in_r_bits_resp; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_in_r_bits_last; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_aw_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_out_aw_bits_addr; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_w_valid; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_out_w_bits_data; // @[Buffer.scala 58:29]
  wire [3:0] axi4buf_12_auto_out_w_bits_strb; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_b_bits_id; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_ar_bits_id; // @[Buffer.scala 58:29]
  wire [29:0] axi4buf_12_auto_out_ar_bits_addr; // @[Buffer.scala 58:29]
  wire [2:0] axi4buf_12_auto_out_ar_bits_size; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_ready; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_valid; // @[Buffer.scala 58:29]
  wire  axi4buf_12_auto_out_r_bits_id; // @[Buffer.scala 58:29]
  wire [31:0] axi4buf_12_auto_out_r_bits_data; // @[Buffer.scala 58:29]
  wire  buffer_clock; // @[Buffer.scala 29:28]
  wire  buffer_reset; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_clock; // @[Buffer.scala 29:28]
  wire  buffer_1_reset; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_1_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_1_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_1_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_clock; // @[Buffer.scala 29:28]
  wire  buffer_2_reset; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_2_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_2_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_clock; // @[Buffer.scala 29:28]
  wire  buffer_3_reset; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_3_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_3_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_3_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_4_clock; // @[Buffer.scala 29:28]
  wire  buffer_4_reset; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_4_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_4_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_4_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_5_clock; // @[Buffer.scala 29:28]
  wire  buffer_5_reset; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_5_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_5_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_5_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_6_clock; // @[Buffer.scala 29:28]
  wire  buffer_6_reset; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_6_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_6_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_6_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_7_clock; // @[Buffer.scala 29:28]
  wire  buffer_7_reset; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_7_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_7_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_7_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_8_clock; // @[Buffer.scala 29:28]
  wire  buffer_8_reset; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_8_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_8_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_8_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_9_clock; // @[Buffer.scala 29:28]
  wire  buffer_9_reset; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_9_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_9_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_9_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_10_clock; // @[Buffer.scala 29:28]
  wire  buffer_10_reset; // @[Buffer.scala 29:28]
  wire  buffer_10_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_10_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_10_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_10_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_10_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_10_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_10_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_10_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_11_clock; // @[Buffer.scala 29:28]
  wire  buffer_11_reset; // @[Buffer.scala 29:28]
  wire  buffer_11_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_11_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_11_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_11_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_11_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_11_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_11_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_11_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_12_clock; // @[Buffer.scala 29:28]
  wire  buffer_12_reset; // @[Buffer.scala 29:28]
  wire  buffer_12_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_12_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_12_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_12_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_12_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_12_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_12_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_12_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_13_clock; // @[Buffer.scala 29:28]
  wire  buffer_13_reset; // @[Buffer.scala 29:28]
  wire  buffer_13_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_13_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_13_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_13_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_13_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_13_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_13_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_13_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_14_clock; // @[Buffer.scala 29:28]
  wire  buffer_14_reset; // @[Buffer.scala 29:28]
  wire  buffer_14_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_14_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_14_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_14_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_14_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_14_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_14_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_14_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_15_clock; // @[Buffer.scala 29:28]
  wire  buffer_15_reset; // @[Buffer.scala 29:28]
  wire  buffer_15_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_15_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_15_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_15_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_15_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_15_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_15_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_15_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_16_clock; // @[Buffer.scala 29:28]
  wire  buffer_16_reset; // @[Buffer.scala 29:28]
  wire  buffer_16_auto_in_ready; // @[Buffer.scala 29:28]
  wire  buffer_16_auto_in_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_16_auto_in_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_16_auto_in_bits_last; // @[Buffer.scala 29:28]
  wire  buffer_16_auto_out_ready; // @[Buffer.scala 29:28]
  wire  buffer_16_auto_out_valid; // @[Buffer.scala 29:28]
  wire [31:0] buffer_16_auto_out_bits_data; // @[Buffer.scala 29:28]
  wire  buffer_16_auto_out_bits_last; // @[Buffer.scala 29:28]
  wire  converter_auto_in_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_aw_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_aw_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_aw_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_in_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_in_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_in_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_in_ar_bits_id; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_in_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_in_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_in_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_in_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_in_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_in_r_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_aw_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_aw_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_aw_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_w_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_w_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_w_bits_data; // @[Node.scala 65:31]
  wire [3:0] converter_auto_out_w_bits_strb; // @[Node.scala 65:31]
  wire  converter_auto_out_w_bits_last; // @[Node.scala 65:31]
  wire  converter_auto_out_b_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_b_valid; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_b_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_valid; // @[Node.scala 65:31]
  wire  converter_auto_out_ar_bits_id; // @[Node.scala 65:31]
  wire [29:0] converter_auto_out_ar_bits_addr; // @[Node.scala 65:31]
  wire [2:0] converter_auto_out_ar_bits_size; // @[Node.scala 65:31]
  wire  converter_auto_out_r_ready; // @[Node.scala 65:31]
  wire  converter_auto_out_r_valid; // @[Node.scala 65:31]
  wire [31:0] converter_auto_out_r_bits_data; // @[Node.scala 65:31]
  wire [1:0] converter_auto_out_r_bits_resp; // @[Node.scala 65:31]
  wire  converter_auto_out_r_bits_last; // @[Node.scala 65:31]
  wire  converter_1_auto_in_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_valid; // @[Nodes.scala 165:31]
  wire [7:0] converter_1_auto_in_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_in_bits_last; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_ready; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_valid; // @[Nodes.scala 165:31]
  wire [7:0] converter_1_auto_out_bits_data; // @[Nodes.scala 165:31]
  wire  converter_1_auto_out_bits_last; // @[Nodes.scala 165:31]
  wire  converter_2_auto_in_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_in_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_in_bits_last; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_ready; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_valid; // @[Nodes.scala 201:31]
  wire [7:0] converter_2_auto_out_bits_data; // @[Nodes.scala 201:31]
  wire  converter_2_auto_out_bits_last; // @[Nodes.scala 201:31]
  wire  converter_3_auto_in_ready; // @[Nodes.scala 165:31]
  wire  converter_3_auto_in_valid; // @[Nodes.scala 165:31]
  wire [31:0] converter_3_auto_in_bits_data; // @[Nodes.scala 165:31]
  wire  converter_3_auto_in_bits_last; // @[Nodes.scala 165:31]
  wire  converter_3_auto_out_ready; // @[Nodes.scala 165:31]
  wire  converter_3_auto_out_valid; // @[Nodes.scala 165:31]
  wire [31:0] converter_3_auto_out_bits_data; // @[Nodes.scala 165:31]
  wire  converter_3_auto_out_bits_last; // @[Nodes.scala 165:31]
  wire  converter_4_auto_in_ready; // @[Nodes.scala 165:31]
  wire  converter_4_auto_in_valid; // @[Nodes.scala 165:31]
  wire [31:0] converter_4_auto_in_bits_data; // @[Nodes.scala 165:31]
  wire  converter_4_auto_in_bits_last; // @[Nodes.scala 165:31]
  wire  converter_4_auto_out_ready; // @[Nodes.scala 165:31]
  wire  converter_4_auto_out_valid; // @[Nodes.scala 165:31]
  wire [31:0] converter_4_auto_out_bits_data; // @[Nodes.scala 165:31]
  wire  converter_4_auto_out_bits_last; // @[Nodes.scala 165:31]
  AXI4StreamWidthAdapater_4_to_1 widthAdapter ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_clock),
    .reset(widthAdapter_reset),
    .auto_in_ready(widthAdapter_auto_in_ready),
    .auto_in_valid(widthAdapter_auto_in_valid),
    .auto_in_bits_data(widthAdapter_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_auto_in_bits_last),
    .auto_out_ready(widthAdapter_auto_out_ready),
    .auto_out_valid(widthAdapter_auto_out_valid),
    .auto_out_bits_data(widthAdapter_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_auto_out_bits_last)
  );
  AXI4Splitter in_split ( // @[LISTestWithLA.scala 55:29]
    .clock(in_split_clock),
    .reset(in_split_reset),
    .auto_mem_in_aw_ready(in_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(in_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(in_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(in_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(in_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(in_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(in_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(in_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(in_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(in_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(in_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(in_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(in_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(in_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(in_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(in_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(in_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(in_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(in_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(in_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(in_split_auto_stream_in_ready),
    .auto_stream_in_valid(in_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(in_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(in_split_auto_stream_in_bits_last),
    .auto_stream_out_4_ready(in_split_auto_stream_out_4_ready),
    .auto_stream_out_4_valid(in_split_auto_stream_out_4_valid),
    .auto_stream_out_4_bits_data(in_split_auto_stream_out_4_bits_data),
    .auto_stream_out_4_bits_last(in_split_auto_stream_out_4_bits_last),
    .auto_stream_out_3_ready(in_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(in_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(in_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(in_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(in_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(in_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(in_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(in_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(in_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(in_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(in_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(in_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(in_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(in_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(in_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(in_split_auto_stream_out_0_bits_last)
  );
  StreamBuffer in_queue ( // @[LISTestWithLA.scala 56:29]
    .clock(in_queue_clock),
    .reset(in_queue_reset),
    .auto_out_out_ready(in_queue_auto_out_out_ready),
    .auto_out_out_valid(in_queue_auto_out_out_valid),
    .auto_out_out_bits_data(in_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(in_queue_auto_out_out_bits_last),
    .auto_in_in_ready(in_queue_auto_in_in_ready),
    .auto_in_in_valid(in_queue_auto_in_in_valid),
    .auto_in_in_bits_data(in_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(in_queue_auto_in_in_bits_last)
  );
  AXI4LISBlock lisFifo ( // @[LISTestWithLA.scala 59:33]
    .clock(lisFifo_clock),
    .reset(lisFifo_reset),
    .auto_mem_in_aw_ready(lisFifo_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(lisFifo_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(lisFifo_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(lisFifo_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(lisFifo_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(lisFifo_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(lisFifo_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(lisFifo_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(lisFifo_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(lisFifo_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(lisFifo_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(lisFifo_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(lisFifo_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(lisFifo_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(lisFifo_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(lisFifo_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(lisFifo_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(lisFifo_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(lisFifo_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(lisFifo_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(lisFifo_auto_stream_in_ready),
    .auto_stream_in_valid(lisFifo_auto_stream_in_valid),
    .auto_stream_in_bits_data(lisFifo_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(lisFifo_auto_stream_in_bits_last),
    .auto_stream_out_ready(lisFifo_auto_stream_out_ready),
    .auto_stream_out_valid(lisFifo_auto_stream_out_valid),
    .auto_stream_out_bits_data(lisFifo_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(lisFifo_auto_stream_out_bits_last)
  );
  AXI4StreamMux lisFifo_mux0 ( // @[LISTestWithLA.scala 60:33]
    .clock(lisFifo_mux0_clock),
    .reset(lisFifo_mux0_reset),
    .auto_register_in_aw_ready(lisFifo_mux0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(lisFifo_mux0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(lisFifo_mux0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(lisFifo_mux0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(lisFifo_mux0_auto_register_in_w_ready),
    .auto_register_in_w_valid(lisFifo_mux0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(lisFifo_mux0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(lisFifo_mux0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(lisFifo_mux0_auto_register_in_b_ready),
    .auto_register_in_b_valid(lisFifo_mux0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(lisFifo_mux0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(lisFifo_mux0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(lisFifo_mux0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(lisFifo_mux0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(lisFifo_mux0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(lisFifo_mux0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(lisFifo_mux0_auto_register_in_r_ready),
    .auto_register_in_r_valid(lisFifo_mux0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(lisFifo_mux0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(lisFifo_mux0_auto_register_in_r_bits_data),
    .auto_stream_in_4_ready(lisFifo_mux0_auto_stream_in_4_ready),
    .auto_stream_in_4_valid(lisFifo_mux0_auto_stream_in_4_valid),
    .auto_stream_in_4_bits_data(lisFifo_mux0_auto_stream_in_4_bits_data),
    .auto_stream_in_4_bits_last(lisFifo_mux0_auto_stream_in_4_bits_last),
    .auto_stream_in_3_ready(lisFifo_mux0_auto_stream_in_3_ready),
    .auto_stream_in_3_valid(lisFifo_mux0_auto_stream_in_3_valid),
    .auto_stream_in_3_bits_data(lisFifo_mux0_auto_stream_in_3_bits_data),
    .auto_stream_in_3_bits_last(lisFifo_mux0_auto_stream_in_3_bits_last),
    .auto_stream_in_2_ready(lisFifo_mux0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(lisFifo_mux0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(lisFifo_mux0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(lisFifo_mux0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(lisFifo_mux0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(lisFifo_mux0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(lisFifo_mux0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(lisFifo_mux0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(lisFifo_mux0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(lisFifo_mux0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(lisFifo_mux0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(lisFifo_mux0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(lisFifo_mux0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(lisFifo_mux0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(lisFifo_mux0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(lisFifo_mux0_auto_stream_out_0_bits_last)
  );
  AXI4LISBlock_1 lisInput ( // @[LISTestWithLA.scala 66:34]
    .clock(lisInput_clock),
    .reset(lisInput_reset),
    .auto_mem_in_aw_ready(lisInput_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(lisInput_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(lisInput_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(lisInput_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(lisInput_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(lisInput_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(lisInput_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(lisInput_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(lisInput_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(lisInput_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(lisInput_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(lisInput_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(lisInput_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(lisInput_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(lisInput_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(lisInput_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(lisInput_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(lisInput_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(lisInput_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(lisInput_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(lisInput_auto_stream_in_ready),
    .auto_stream_in_valid(lisInput_auto_stream_in_valid),
    .auto_stream_in_bits_data(lisInput_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(lisInput_auto_stream_in_bits_last),
    .auto_stream_out_ready(lisInput_auto_stream_out_ready),
    .auto_stream_out_valid(lisInput_auto_stream_out_valid),
    .auto_stream_out_bits_data(lisInput_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(lisInput_auto_stream_out_bits_last)
  );
  AXI4StreamMux lisInput_mux0 ( // @[LISTestWithLA.scala 67:34]
    .clock(lisInput_mux0_clock),
    .reset(lisInput_mux0_reset),
    .auto_register_in_aw_ready(lisInput_mux0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(lisInput_mux0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(lisInput_mux0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(lisInput_mux0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(lisInput_mux0_auto_register_in_w_ready),
    .auto_register_in_w_valid(lisInput_mux0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(lisInput_mux0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(lisInput_mux0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(lisInput_mux0_auto_register_in_b_ready),
    .auto_register_in_b_valid(lisInput_mux0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(lisInput_mux0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(lisInput_mux0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(lisInput_mux0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(lisInput_mux0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(lisInput_mux0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(lisInput_mux0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(lisInput_mux0_auto_register_in_r_ready),
    .auto_register_in_r_valid(lisInput_mux0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(lisInput_mux0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(lisInput_mux0_auto_register_in_r_bits_data),
    .auto_stream_in_4_ready(lisInput_mux0_auto_stream_in_4_ready),
    .auto_stream_in_4_valid(lisInput_mux0_auto_stream_in_4_valid),
    .auto_stream_in_4_bits_data(lisInput_mux0_auto_stream_in_4_bits_data),
    .auto_stream_in_4_bits_last(lisInput_mux0_auto_stream_in_4_bits_last),
    .auto_stream_in_3_ready(lisInput_mux0_auto_stream_in_3_ready),
    .auto_stream_in_3_valid(lisInput_mux0_auto_stream_in_3_valid),
    .auto_stream_in_3_bits_data(lisInput_mux0_auto_stream_in_3_bits_data),
    .auto_stream_in_3_bits_last(lisInput_mux0_auto_stream_in_3_bits_last),
    .auto_stream_in_2_ready(lisInput_mux0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(lisInput_mux0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(lisInput_mux0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(lisInput_mux0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(lisInput_mux0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(lisInput_mux0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(lisInput_mux0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(lisInput_mux0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(lisInput_mux0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(lisInput_mux0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(lisInput_mux0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(lisInput_mux0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(lisInput_mux0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(lisInput_mux0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(lisInput_mux0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(lisInput_mux0_auto_stream_out_0_bits_last)
  );
  AXI4LISBlock_2 lisFixed ( // @[LISTestWithLA.scala 73:34]
    .clock(lisFixed_clock),
    .reset(lisFixed_reset),
    .auto_mem_in_aw_ready(lisFixed_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(lisFixed_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(lisFixed_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(lisFixed_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(lisFixed_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(lisFixed_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(lisFixed_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(lisFixed_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(lisFixed_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(lisFixed_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(lisFixed_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(lisFixed_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(lisFixed_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(lisFixed_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(lisFixed_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(lisFixed_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(lisFixed_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(lisFixed_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(lisFixed_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(lisFixed_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(lisFixed_auto_stream_in_ready),
    .auto_stream_in_valid(lisFixed_auto_stream_in_valid),
    .auto_stream_in_bits_data(lisFixed_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(lisFixed_auto_stream_in_bits_last),
    .auto_stream_out_ready(lisFixed_auto_stream_out_ready),
    .auto_stream_out_valid(lisFixed_auto_stream_out_valid),
    .auto_stream_out_bits_data(lisFixed_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(lisFixed_auto_stream_out_bits_last)
  );
  AXI4StreamMux lisFixed_mux0 ( // @[LISTestWithLA.scala 74:34]
    .clock(lisFixed_mux0_clock),
    .reset(lisFixed_mux0_reset),
    .auto_register_in_aw_ready(lisFixed_mux0_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(lisFixed_mux0_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(lisFixed_mux0_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(lisFixed_mux0_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(lisFixed_mux0_auto_register_in_w_ready),
    .auto_register_in_w_valid(lisFixed_mux0_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(lisFixed_mux0_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(lisFixed_mux0_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(lisFixed_mux0_auto_register_in_b_ready),
    .auto_register_in_b_valid(lisFixed_mux0_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(lisFixed_mux0_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(lisFixed_mux0_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(lisFixed_mux0_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(lisFixed_mux0_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(lisFixed_mux0_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(lisFixed_mux0_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(lisFixed_mux0_auto_register_in_r_ready),
    .auto_register_in_r_valid(lisFixed_mux0_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(lisFixed_mux0_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(lisFixed_mux0_auto_register_in_r_bits_data),
    .auto_stream_in_4_ready(lisFixed_mux0_auto_stream_in_4_ready),
    .auto_stream_in_4_valid(lisFixed_mux0_auto_stream_in_4_valid),
    .auto_stream_in_4_bits_data(lisFixed_mux0_auto_stream_in_4_bits_data),
    .auto_stream_in_4_bits_last(lisFixed_mux0_auto_stream_in_4_bits_last),
    .auto_stream_in_3_ready(lisFixed_mux0_auto_stream_in_3_ready),
    .auto_stream_in_3_valid(lisFixed_mux0_auto_stream_in_3_valid),
    .auto_stream_in_3_bits_data(lisFixed_mux0_auto_stream_in_3_bits_data),
    .auto_stream_in_3_bits_last(lisFixed_mux0_auto_stream_in_3_bits_last),
    .auto_stream_in_2_ready(lisFixed_mux0_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(lisFixed_mux0_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(lisFixed_mux0_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(lisFixed_mux0_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(lisFixed_mux0_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(lisFixed_mux0_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(lisFixed_mux0_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(lisFixed_mux0_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(lisFixed_mux0_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(lisFixed_mux0_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(lisFixed_mux0_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(lisFixed_mux0_auto_stream_in_0_bits_last),
    .auto_stream_out_0_ready(lisFixed_mux0_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(lisFixed_mux0_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(lisFixed_mux0_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(lisFixed_mux0_auto_stream_out_0_bits_last)
  );
  AXI4StreamBIST bist ( // @[LISTestWithLA.scala 79:34]
    .clock(bist_clock),
    .reset(bist_reset),
    .auto_mem_in_aw_ready(bist_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(bist_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(bist_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(bist_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(bist_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(bist_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(bist_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(bist_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(bist_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(bist_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(bist_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(bist_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(bist_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(bist_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(bist_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(bist_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(bist_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(bist_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(bist_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(bist_auto_mem_in_r_bits_data),
    .auto_stream_out_ready(bist_auto_stream_out_ready),
    .auto_stream_out_valid(bist_auto_stream_out_valid),
    .auto_stream_out_bits_data(bist_auto_stream_out_bits_data),
    .auto_stream_out_bits_last(bist_auto_stream_out_bits_last)
  );
  AXI4Splitter_1 bist_split ( // @[LISTestWithLA.scala 80:34]
    .clock(bist_split_clock),
    .reset(bist_split_reset),
    .auto_mem_in_aw_ready(bist_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(bist_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(bist_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(bist_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(bist_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(bist_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(bist_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(bist_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(bist_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(bist_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(bist_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(bist_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(bist_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(bist_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(bist_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(bist_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(bist_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(bist_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(bist_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(bist_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(bist_split_auto_stream_in_ready),
    .auto_stream_in_valid(bist_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(bist_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(bist_split_auto_stream_in_bits_last),
    .auto_stream_out_3_ready(bist_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(bist_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(bist_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(bist_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(bist_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(bist_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(bist_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(bist_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(bist_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(bist_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(bist_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(bist_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(bist_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(bist_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(bist_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(bist_split_auto_stream_out_0_bits_last)
  );
  AXI4StreamMux_3 out_mux ( // @[LISTestWithLA.scala 83:29]
    .clock(out_mux_clock),
    .reset(out_mux_reset),
    .auto_register_in_aw_ready(out_mux_auto_register_in_aw_ready),
    .auto_register_in_aw_valid(out_mux_auto_register_in_aw_valid),
    .auto_register_in_aw_bits_id(out_mux_auto_register_in_aw_bits_id),
    .auto_register_in_aw_bits_addr(out_mux_auto_register_in_aw_bits_addr),
    .auto_register_in_w_ready(out_mux_auto_register_in_w_ready),
    .auto_register_in_w_valid(out_mux_auto_register_in_w_valid),
    .auto_register_in_w_bits_data(out_mux_auto_register_in_w_bits_data),
    .auto_register_in_w_bits_strb(out_mux_auto_register_in_w_bits_strb),
    .auto_register_in_b_ready(out_mux_auto_register_in_b_ready),
    .auto_register_in_b_valid(out_mux_auto_register_in_b_valid),
    .auto_register_in_b_bits_id(out_mux_auto_register_in_b_bits_id),
    .auto_register_in_ar_ready(out_mux_auto_register_in_ar_ready),
    .auto_register_in_ar_valid(out_mux_auto_register_in_ar_valid),
    .auto_register_in_ar_bits_id(out_mux_auto_register_in_ar_bits_id),
    .auto_register_in_ar_bits_addr(out_mux_auto_register_in_ar_bits_addr),
    .auto_register_in_ar_bits_size(out_mux_auto_register_in_ar_bits_size),
    .auto_register_in_r_ready(out_mux_auto_register_in_r_ready),
    .auto_register_in_r_valid(out_mux_auto_register_in_r_valid),
    .auto_register_in_r_bits_id(out_mux_auto_register_in_r_bits_id),
    .auto_register_in_r_bits_data(out_mux_auto_register_in_r_bits_data),
    .auto_stream_in_5_ready(out_mux_auto_stream_in_5_ready),
    .auto_stream_in_5_valid(out_mux_auto_stream_in_5_valid),
    .auto_stream_in_5_bits_data(out_mux_auto_stream_in_5_bits_data),
    .auto_stream_in_5_bits_last(out_mux_auto_stream_in_5_bits_last),
    .auto_stream_in_4_ready(out_mux_auto_stream_in_4_ready),
    .auto_stream_in_4_valid(out_mux_auto_stream_in_4_valid),
    .auto_stream_in_4_bits_data(out_mux_auto_stream_in_4_bits_data),
    .auto_stream_in_4_bits_last(out_mux_auto_stream_in_4_bits_last),
    .auto_stream_in_3_ready(out_mux_auto_stream_in_3_ready),
    .auto_stream_in_3_valid(out_mux_auto_stream_in_3_valid),
    .auto_stream_in_3_bits_data(out_mux_auto_stream_in_3_bits_data),
    .auto_stream_in_3_bits_last(out_mux_auto_stream_in_3_bits_last),
    .auto_stream_in_2_ready(out_mux_auto_stream_in_2_ready),
    .auto_stream_in_2_valid(out_mux_auto_stream_in_2_valid),
    .auto_stream_in_2_bits_data(out_mux_auto_stream_in_2_bits_data),
    .auto_stream_in_2_bits_last(out_mux_auto_stream_in_2_bits_last),
    .auto_stream_in_1_ready(out_mux_auto_stream_in_1_ready),
    .auto_stream_in_1_valid(out_mux_auto_stream_in_1_valid),
    .auto_stream_in_1_bits_data(out_mux_auto_stream_in_1_bits_data),
    .auto_stream_in_1_bits_last(out_mux_auto_stream_in_1_bits_last),
    .auto_stream_in_0_ready(out_mux_auto_stream_in_0_ready),
    .auto_stream_in_0_valid(out_mux_auto_stream_in_0_valid),
    .auto_stream_in_0_bits_data(out_mux_auto_stream_in_0_bits_data),
    .auto_stream_in_0_bits_last(out_mux_auto_stream_in_0_bits_last),
    .auto_stream_out_1_ready(out_mux_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(out_mux_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(out_mux_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(out_mux_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(out_mux_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(out_mux_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(out_mux_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(out_mux_auto_stream_out_0_bits_last)
  );
  AXI4Splitter_2 out_split ( // @[LISTestWithLA.scala 84:29]
    .clock(out_split_clock),
    .reset(out_split_reset),
    .auto_mem_in_aw_ready(out_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(out_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(out_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(out_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(out_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(out_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(out_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(out_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(out_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(out_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(out_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(out_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(out_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(out_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(out_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(out_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(out_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(out_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(out_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(out_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(out_split_auto_stream_in_ready),
    .auto_stream_in_valid(out_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(out_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(out_split_auto_stream_in_bits_last),
    .auto_stream_out_1_ready(out_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(out_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(out_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(out_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(out_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(out_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(out_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(out_split_auto_stream_out_0_bits_last)
  );
  StreamBuffer_1 out_queue ( // @[LISTestWithLA.scala 85:29]
    .clock(out_queue_clock),
    .reset(out_queue_reset),
    .auto_out_out_ready(out_queue_auto_out_out_ready),
    .auto_out_out_valid(out_queue_auto_out_out_valid),
    .auto_out_out_bits_data(out_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(out_queue_auto_out_out_bits_last),
    .auto_in_in_ready(out_queue_auto_in_in_ready),
    .auto_in_in_valid(out_queue_auto_in_in_valid),
    .auto_in_in_bits_data(out_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(out_queue_auto_in_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_4 widthAdapter_1 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_1_clock),
    .reset(widthAdapter_1_reset),
    .auto_in_ready(widthAdapter_1_auto_in_ready),
    .auto_in_valid(widthAdapter_1_auto_in_valid),
    .auto_in_bits_data(widthAdapter_1_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_1_auto_in_bits_last),
    .auto_out_ready(widthAdapter_1_auto_out_ready),
    .auto_out_valid(widthAdapter_1_auto_out_valid),
    .auto_out_bits_data(widthAdapter_1_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_1_auto_out_bits_last)
  );
  StreamBuffer_2 uTx_queue ( // @[LISTestWithLA.scala 89:29]
    .clock(uTx_queue_clock),
    .reset(uTx_queue_reset),
    .auto_out_out_ready(uTx_queue_auto_out_out_ready),
    .auto_out_out_valid(uTx_queue_auto_out_out_valid),
    .auto_out_out_bits_data(uTx_queue_auto_out_out_bits_data),
    .auto_out_out_bits_last(uTx_queue_auto_out_out_bits_last),
    .auto_in_in_ready(uTx_queue_auto_in_in_ready),
    .auto_in_in_valid(uTx_queue_auto_in_in_valid),
    .auto_in_in_bits_data(uTx_queue_auto_in_in_bits_data),
    .auto_in_in_bits_last(uTx_queue_auto_in_in_bits_last)
  );
  AXI4StreamWidthAdapater_1_to_4 widthAdapter_2 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_2_clock),
    .reset(widthAdapter_2_reset),
    .auto_in_ready(widthAdapter_2_auto_in_ready),
    .auto_in_valid(widthAdapter_2_auto_in_valid),
    .auto_in_bits_data(widthAdapter_2_auto_in_bits_data),
    .auto_in_bits_last(widthAdapter_2_auto_in_bits_last),
    .auto_out_ready(widthAdapter_2_auto_out_ready),
    .auto_out_valid(widthAdapter_2_auto_out_valid),
    .auto_out_bits_data(widthAdapter_2_auto_out_bits_data),
    .auto_out_bits_last(widthAdapter_2_auto_out_bits_last)
  );
  AXI4StreamWidthAdapater_4_to_1_1 widthAdapter_3 ( // @[AXI4StreamWidthAdapter.scala 82:34]
    .clock(widthAdapter_3_clock),
    .reset(widthAdapter_3_reset),
    .auto_in_ready(widthAdapter_3_auto_in_ready),
    .auto_in_valid(widthAdapter_3_auto_in_valid),
    .auto_in_bits_data(widthAdapter_3_auto_in_bits_data),
    .auto_out_ready(widthAdapter_3_auto_out_ready),
    .auto_out_valid(widthAdapter_3_auto_out_valid),
    .auto_out_bits_data(widthAdapter_3_auto_out_bits_data)
  );
  AXI4Splitter_1 uRx_split ( // @[LISTestWithLA.scala 92:29]
    .clock(uRx_split_clock),
    .reset(uRx_split_reset),
    .auto_mem_in_aw_ready(uRx_split_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(uRx_split_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(uRx_split_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(uRx_split_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(uRx_split_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(uRx_split_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(uRx_split_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(uRx_split_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(uRx_split_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(uRx_split_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(uRx_split_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(uRx_split_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(uRx_split_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(uRx_split_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(uRx_split_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(uRx_split_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(uRx_split_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(uRx_split_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(uRx_split_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(uRx_split_auto_mem_in_r_bits_data),
    .auto_stream_in_ready(uRx_split_auto_stream_in_ready),
    .auto_stream_in_valid(uRx_split_auto_stream_in_valid),
    .auto_stream_in_bits_data(uRx_split_auto_stream_in_bits_data),
    .auto_stream_in_bits_last(uRx_split_auto_stream_in_bits_last),
    .auto_stream_out_3_ready(uRx_split_auto_stream_out_3_ready),
    .auto_stream_out_3_valid(uRx_split_auto_stream_out_3_valid),
    .auto_stream_out_3_bits_data(uRx_split_auto_stream_out_3_bits_data),
    .auto_stream_out_3_bits_last(uRx_split_auto_stream_out_3_bits_last),
    .auto_stream_out_2_ready(uRx_split_auto_stream_out_2_ready),
    .auto_stream_out_2_valid(uRx_split_auto_stream_out_2_valid),
    .auto_stream_out_2_bits_data(uRx_split_auto_stream_out_2_bits_data),
    .auto_stream_out_2_bits_last(uRx_split_auto_stream_out_2_bits_last),
    .auto_stream_out_1_ready(uRx_split_auto_stream_out_1_ready),
    .auto_stream_out_1_valid(uRx_split_auto_stream_out_1_valid),
    .auto_stream_out_1_bits_data(uRx_split_auto_stream_out_1_bits_data),
    .auto_stream_out_1_bits_last(uRx_split_auto_stream_out_1_bits_last),
    .auto_stream_out_0_ready(uRx_split_auto_stream_out_0_ready),
    .auto_stream_out_0_valid(uRx_split_auto_stream_out_0_valid),
    .auto_stream_out_0_bits_data(uRx_split_auto_stream_out_0_bits_data),
    .auto_stream_out_0_bits_last(uRx_split_auto_stream_out_0_bits_last)
  );
  AXI4UARTBlock uart ( // @[LISTestWithLA.scala 93:29]
    .clock(uart_clock),
    .reset(uart_reset),
    .auto_mem_in_aw_ready(uart_auto_mem_in_aw_ready),
    .auto_mem_in_aw_valid(uart_auto_mem_in_aw_valid),
    .auto_mem_in_aw_bits_id(uart_auto_mem_in_aw_bits_id),
    .auto_mem_in_aw_bits_addr(uart_auto_mem_in_aw_bits_addr),
    .auto_mem_in_w_ready(uart_auto_mem_in_w_ready),
    .auto_mem_in_w_valid(uart_auto_mem_in_w_valid),
    .auto_mem_in_w_bits_data(uart_auto_mem_in_w_bits_data),
    .auto_mem_in_w_bits_strb(uart_auto_mem_in_w_bits_strb),
    .auto_mem_in_b_ready(uart_auto_mem_in_b_ready),
    .auto_mem_in_b_valid(uart_auto_mem_in_b_valid),
    .auto_mem_in_b_bits_id(uart_auto_mem_in_b_bits_id),
    .auto_mem_in_ar_ready(uart_auto_mem_in_ar_ready),
    .auto_mem_in_ar_valid(uart_auto_mem_in_ar_valid),
    .auto_mem_in_ar_bits_id(uart_auto_mem_in_ar_bits_id),
    .auto_mem_in_ar_bits_addr(uart_auto_mem_in_ar_bits_addr),
    .auto_mem_in_ar_bits_size(uart_auto_mem_in_ar_bits_size),
    .auto_mem_in_r_ready(uart_auto_mem_in_r_ready),
    .auto_mem_in_r_valid(uart_auto_mem_in_r_valid),
    .auto_mem_in_r_bits_id(uart_auto_mem_in_r_bits_id),
    .auto_mem_in_r_bits_data(uart_auto_mem_in_r_bits_data),
    .auto_in_in_ready(uart_auto_in_in_ready),
    .auto_in_in_valid(uart_auto_in_in_valid),
    .auto_in_in_bits_data(uart_auto_in_in_bits_data),
    .auto_out_out_ready(uart_auto_out_out_ready),
    .auto_out_out_valid(uart_auto_out_out_valid),
    .auto_out_out_bits_data(uart_auto_out_out_bits_data),
    .int_0(uart_int_0),
    .io_txd(uart_io_txd),
    .io_rxd(uart_io_rxd)
  );
  AXI4Xbar bus ( // @[LISTestWithLA.scala 108:23]
    .clock(bus_clock),
    .reset(bus_reset),
    .auto_in_aw_ready(bus_auto_in_aw_ready),
    .auto_in_aw_valid(bus_auto_in_aw_valid),
    .auto_in_aw_bits_id(bus_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(bus_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(bus_auto_in_aw_bits_size),
    .auto_in_w_ready(bus_auto_in_w_ready),
    .auto_in_w_valid(bus_auto_in_w_valid),
    .auto_in_w_bits_data(bus_auto_in_w_bits_data),
    .auto_in_w_bits_strb(bus_auto_in_w_bits_strb),
    .auto_in_w_bits_last(bus_auto_in_w_bits_last),
    .auto_in_b_ready(bus_auto_in_b_ready),
    .auto_in_b_valid(bus_auto_in_b_valid),
    .auto_in_b_bits_resp(bus_auto_in_b_bits_resp),
    .auto_in_ar_ready(bus_auto_in_ar_ready),
    .auto_in_ar_valid(bus_auto_in_ar_valid),
    .auto_in_ar_bits_id(bus_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(bus_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(bus_auto_in_ar_bits_size),
    .auto_in_r_ready(bus_auto_in_r_ready),
    .auto_in_r_valid(bus_auto_in_r_valid),
    .auto_in_r_bits_data(bus_auto_in_r_bits_data),
    .auto_in_r_bits_resp(bus_auto_in_r_bits_resp),
    .auto_in_r_bits_last(bus_auto_in_r_bits_last),
    .auto_out_12_aw_ready(bus_auto_out_12_aw_ready),
    .auto_out_12_aw_valid(bus_auto_out_12_aw_valid),
    .auto_out_12_aw_bits_id(bus_auto_out_12_aw_bits_id),
    .auto_out_12_aw_bits_addr(bus_auto_out_12_aw_bits_addr),
    .auto_out_12_aw_bits_size(bus_auto_out_12_aw_bits_size),
    .auto_out_12_w_ready(bus_auto_out_12_w_ready),
    .auto_out_12_w_valid(bus_auto_out_12_w_valid),
    .auto_out_12_w_bits_data(bus_auto_out_12_w_bits_data),
    .auto_out_12_w_bits_strb(bus_auto_out_12_w_bits_strb),
    .auto_out_12_b_ready(bus_auto_out_12_b_ready),
    .auto_out_12_b_valid(bus_auto_out_12_b_valid),
    .auto_out_12_b_bits_id(bus_auto_out_12_b_bits_id),
    .auto_out_12_b_bits_resp(bus_auto_out_12_b_bits_resp),
    .auto_out_12_ar_ready(bus_auto_out_12_ar_ready),
    .auto_out_12_ar_valid(bus_auto_out_12_ar_valid),
    .auto_out_12_ar_bits_id(bus_auto_out_12_ar_bits_id),
    .auto_out_12_ar_bits_addr(bus_auto_out_12_ar_bits_addr),
    .auto_out_12_ar_bits_size(bus_auto_out_12_ar_bits_size),
    .auto_out_12_r_ready(bus_auto_out_12_r_ready),
    .auto_out_12_r_valid(bus_auto_out_12_r_valid),
    .auto_out_12_r_bits_id(bus_auto_out_12_r_bits_id),
    .auto_out_12_r_bits_data(bus_auto_out_12_r_bits_data),
    .auto_out_12_r_bits_resp(bus_auto_out_12_r_bits_resp),
    .auto_out_12_r_bits_last(bus_auto_out_12_r_bits_last),
    .auto_out_11_aw_ready(bus_auto_out_11_aw_ready),
    .auto_out_11_aw_valid(bus_auto_out_11_aw_valid),
    .auto_out_11_aw_bits_id(bus_auto_out_11_aw_bits_id),
    .auto_out_11_aw_bits_addr(bus_auto_out_11_aw_bits_addr),
    .auto_out_11_aw_bits_size(bus_auto_out_11_aw_bits_size),
    .auto_out_11_w_ready(bus_auto_out_11_w_ready),
    .auto_out_11_w_valid(bus_auto_out_11_w_valid),
    .auto_out_11_w_bits_data(bus_auto_out_11_w_bits_data),
    .auto_out_11_w_bits_strb(bus_auto_out_11_w_bits_strb),
    .auto_out_11_b_ready(bus_auto_out_11_b_ready),
    .auto_out_11_b_valid(bus_auto_out_11_b_valid),
    .auto_out_11_b_bits_id(bus_auto_out_11_b_bits_id),
    .auto_out_11_b_bits_resp(bus_auto_out_11_b_bits_resp),
    .auto_out_11_ar_ready(bus_auto_out_11_ar_ready),
    .auto_out_11_ar_valid(bus_auto_out_11_ar_valid),
    .auto_out_11_ar_bits_id(bus_auto_out_11_ar_bits_id),
    .auto_out_11_ar_bits_addr(bus_auto_out_11_ar_bits_addr),
    .auto_out_11_ar_bits_size(bus_auto_out_11_ar_bits_size),
    .auto_out_11_r_ready(bus_auto_out_11_r_ready),
    .auto_out_11_r_valid(bus_auto_out_11_r_valid),
    .auto_out_11_r_bits_id(bus_auto_out_11_r_bits_id),
    .auto_out_11_r_bits_data(bus_auto_out_11_r_bits_data),
    .auto_out_11_r_bits_resp(bus_auto_out_11_r_bits_resp),
    .auto_out_11_r_bits_last(bus_auto_out_11_r_bits_last),
    .auto_out_10_aw_ready(bus_auto_out_10_aw_ready),
    .auto_out_10_aw_valid(bus_auto_out_10_aw_valid),
    .auto_out_10_aw_bits_id(bus_auto_out_10_aw_bits_id),
    .auto_out_10_aw_bits_addr(bus_auto_out_10_aw_bits_addr),
    .auto_out_10_aw_bits_size(bus_auto_out_10_aw_bits_size),
    .auto_out_10_w_ready(bus_auto_out_10_w_ready),
    .auto_out_10_w_valid(bus_auto_out_10_w_valid),
    .auto_out_10_w_bits_data(bus_auto_out_10_w_bits_data),
    .auto_out_10_w_bits_strb(bus_auto_out_10_w_bits_strb),
    .auto_out_10_b_ready(bus_auto_out_10_b_ready),
    .auto_out_10_b_valid(bus_auto_out_10_b_valid),
    .auto_out_10_b_bits_id(bus_auto_out_10_b_bits_id),
    .auto_out_10_b_bits_resp(bus_auto_out_10_b_bits_resp),
    .auto_out_10_ar_ready(bus_auto_out_10_ar_ready),
    .auto_out_10_ar_valid(bus_auto_out_10_ar_valid),
    .auto_out_10_ar_bits_id(bus_auto_out_10_ar_bits_id),
    .auto_out_10_ar_bits_addr(bus_auto_out_10_ar_bits_addr),
    .auto_out_10_ar_bits_size(bus_auto_out_10_ar_bits_size),
    .auto_out_10_r_ready(bus_auto_out_10_r_ready),
    .auto_out_10_r_valid(bus_auto_out_10_r_valid),
    .auto_out_10_r_bits_id(bus_auto_out_10_r_bits_id),
    .auto_out_10_r_bits_data(bus_auto_out_10_r_bits_data),
    .auto_out_10_r_bits_resp(bus_auto_out_10_r_bits_resp),
    .auto_out_10_r_bits_last(bus_auto_out_10_r_bits_last),
    .auto_out_9_aw_ready(bus_auto_out_9_aw_ready),
    .auto_out_9_aw_valid(bus_auto_out_9_aw_valid),
    .auto_out_9_aw_bits_id(bus_auto_out_9_aw_bits_id),
    .auto_out_9_aw_bits_addr(bus_auto_out_9_aw_bits_addr),
    .auto_out_9_aw_bits_size(bus_auto_out_9_aw_bits_size),
    .auto_out_9_w_ready(bus_auto_out_9_w_ready),
    .auto_out_9_w_valid(bus_auto_out_9_w_valid),
    .auto_out_9_w_bits_data(bus_auto_out_9_w_bits_data),
    .auto_out_9_w_bits_strb(bus_auto_out_9_w_bits_strb),
    .auto_out_9_b_ready(bus_auto_out_9_b_ready),
    .auto_out_9_b_valid(bus_auto_out_9_b_valid),
    .auto_out_9_b_bits_id(bus_auto_out_9_b_bits_id),
    .auto_out_9_b_bits_resp(bus_auto_out_9_b_bits_resp),
    .auto_out_9_ar_ready(bus_auto_out_9_ar_ready),
    .auto_out_9_ar_valid(bus_auto_out_9_ar_valid),
    .auto_out_9_ar_bits_id(bus_auto_out_9_ar_bits_id),
    .auto_out_9_ar_bits_addr(bus_auto_out_9_ar_bits_addr),
    .auto_out_9_ar_bits_size(bus_auto_out_9_ar_bits_size),
    .auto_out_9_r_ready(bus_auto_out_9_r_ready),
    .auto_out_9_r_valid(bus_auto_out_9_r_valid),
    .auto_out_9_r_bits_id(bus_auto_out_9_r_bits_id),
    .auto_out_9_r_bits_data(bus_auto_out_9_r_bits_data),
    .auto_out_9_r_bits_resp(bus_auto_out_9_r_bits_resp),
    .auto_out_9_r_bits_last(bus_auto_out_9_r_bits_last),
    .auto_out_8_aw_ready(bus_auto_out_8_aw_ready),
    .auto_out_8_aw_valid(bus_auto_out_8_aw_valid),
    .auto_out_8_aw_bits_id(bus_auto_out_8_aw_bits_id),
    .auto_out_8_aw_bits_addr(bus_auto_out_8_aw_bits_addr),
    .auto_out_8_aw_bits_size(bus_auto_out_8_aw_bits_size),
    .auto_out_8_w_ready(bus_auto_out_8_w_ready),
    .auto_out_8_w_valid(bus_auto_out_8_w_valid),
    .auto_out_8_w_bits_data(bus_auto_out_8_w_bits_data),
    .auto_out_8_w_bits_strb(bus_auto_out_8_w_bits_strb),
    .auto_out_8_b_ready(bus_auto_out_8_b_ready),
    .auto_out_8_b_valid(bus_auto_out_8_b_valid),
    .auto_out_8_b_bits_id(bus_auto_out_8_b_bits_id),
    .auto_out_8_b_bits_resp(bus_auto_out_8_b_bits_resp),
    .auto_out_8_ar_ready(bus_auto_out_8_ar_ready),
    .auto_out_8_ar_valid(bus_auto_out_8_ar_valid),
    .auto_out_8_ar_bits_id(bus_auto_out_8_ar_bits_id),
    .auto_out_8_ar_bits_addr(bus_auto_out_8_ar_bits_addr),
    .auto_out_8_ar_bits_size(bus_auto_out_8_ar_bits_size),
    .auto_out_8_r_ready(bus_auto_out_8_r_ready),
    .auto_out_8_r_valid(bus_auto_out_8_r_valid),
    .auto_out_8_r_bits_id(bus_auto_out_8_r_bits_id),
    .auto_out_8_r_bits_data(bus_auto_out_8_r_bits_data),
    .auto_out_8_r_bits_resp(bus_auto_out_8_r_bits_resp),
    .auto_out_8_r_bits_last(bus_auto_out_8_r_bits_last),
    .auto_out_7_aw_ready(bus_auto_out_7_aw_ready),
    .auto_out_7_aw_valid(bus_auto_out_7_aw_valid),
    .auto_out_7_aw_bits_id(bus_auto_out_7_aw_bits_id),
    .auto_out_7_aw_bits_addr(bus_auto_out_7_aw_bits_addr),
    .auto_out_7_aw_bits_size(bus_auto_out_7_aw_bits_size),
    .auto_out_7_w_ready(bus_auto_out_7_w_ready),
    .auto_out_7_w_valid(bus_auto_out_7_w_valid),
    .auto_out_7_w_bits_data(bus_auto_out_7_w_bits_data),
    .auto_out_7_w_bits_strb(bus_auto_out_7_w_bits_strb),
    .auto_out_7_b_ready(bus_auto_out_7_b_ready),
    .auto_out_7_b_valid(bus_auto_out_7_b_valid),
    .auto_out_7_b_bits_id(bus_auto_out_7_b_bits_id),
    .auto_out_7_b_bits_resp(bus_auto_out_7_b_bits_resp),
    .auto_out_7_ar_ready(bus_auto_out_7_ar_ready),
    .auto_out_7_ar_valid(bus_auto_out_7_ar_valid),
    .auto_out_7_ar_bits_id(bus_auto_out_7_ar_bits_id),
    .auto_out_7_ar_bits_addr(bus_auto_out_7_ar_bits_addr),
    .auto_out_7_ar_bits_size(bus_auto_out_7_ar_bits_size),
    .auto_out_7_r_ready(bus_auto_out_7_r_ready),
    .auto_out_7_r_valid(bus_auto_out_7_r_valid),
    .auto_out_7_r_bits_id(bus_auto_out_7_r_bits_id),
    .auto_out_7_r_bits_data(bus_auto_out_7_r_bits_data),
    .auto_out_7_r_bits_resp(bus_auto_out_7_r_bits_resp),
    .auto_out_7_r_bits_last(bus_auto_out_7_r_bits_last),
    .auto_out_6_aw_ready(bus_auto_out_6_aw_ready),
    .auto_out_6_aw_valid(bus_auto_out_6_aw_valid),
    .auto_out_6_aw_bits_id(bus_auto_out_6_aw_bits_id),
    .auto_out_6_aw_bits_addr(bus_auto_out_6_aw_bits_addr),
    .auto_out_6_aw_bits_size(bus_auto_out_6_aw_bits_size),
    .auto_out_6_w_ready(bus_auto_out_6_w_ready),
    .auto_out_6_w_valid(bus_auto_out_6_w_valid),
    .auto_out_6_w_bits_data(bus_auto_out_6_w_bits_data),
    .auto_out_6_w_bits_strb(bus_auto_out_6_w_bits_strb),
    .auto_out_6_b_ready(bus_auto_out_6_b_ready),
    .auto_out_6_b_valid(bus_auto_out_6_b_valid),
    .auto_out_6_b_bits_id(bus_auto_out_6_b_bits_id),
    .auto_out_6_b_bits_resp(bus_auto_out_6_b_bits_resp),
    .auto_out_6_ar_ready(bus_auto_out_6_ar_ready),
    .auto_out_6_ar_valid(bus_auto_out_6_ar_valid),
    .auto_out_6_ar_bits_id(bus_auto_out_6_ar_bits_id),
    .auto_out_6_ar_bits_addr(bus_auto_out_6_ar_bits_addr),
    .auto_out_6_ar_bits_size(bus_auto_out_6_ar_bits_size),
    .auto_out_6_r_ready(bus_auto_out_6_r_ready),
    .auto_out_6_r_valid(bus_auto_out_6_r_valid),
    .auto_out_6_r_bits_id(bus_auto_out_6_r_bits_id),
    .auto_out_6_r_bits_data(bus_auto_out_6_r_bits_data),
    .auto_out_6_r_bits_resp(bus_auto_out_6_r_bits_resp),
    .auto_out_6_r_bits_last(bus_auto_out_6_r_bits_last),
    .auto_out_5_aw_ready(bus_auto_out_5_aw_ready),
    .auto_out_5_aw_valid(bus_auto_out_5_aw_valid),
    .auto_out_5_aw_bits_id(bus_auto_out_5_aw_bits_id),
    .auto_out_5_aw_bits_addr(bus_auto_out_5_aw_bits_addr),
    .auto_out_5_aw_bits_size(bus_auto_out_5_aw_bits_size),
    .auto_out_5_w_ready(bus_auto_out_5_w_ready),
    .auto_out_5_w_valid(bus_auto_out_5_w_valid),
    .auto_out_5_w_bits_data(bus_auto_out_5_w_bits_data),
    .auto_out_5_w_bits_strb(bus_auto_out_5_w_bits_strb),
    .auto_out_5_b_ready(bus_auto_out_5_b_ready),
    .auto_out_5_b_valid(bus_auto_out_5_b_valid),
    .auto_out_5_b_bits_id(bus_auto_out_5_b_bits_id),
    .auto_out_5_b_bits_resp(bus_auto_out_5_b_bits_resp),
    .auto_out_5_ar_ready(bus_auto_out_5_ar_ready),
    .auto_out_5_ar_valid(bus_auto_out_5_ar_valid),
    .auto_out_5_ar_bits_id(bus_auto_out_5_ar_bits_id),
    .auto_out_5_ar_bits_addr(bus_auto_out_5_ar_bits_addr),
    .auto_out_5_ar_bits_size(bus_auto_out_5_ar_bits_size),
    .auto_out_5_r_ready(bus_auto_out_5_r_ready),
    .auto_out_5_r_valid(bus_auto_out_5_r_valid),
    .auto_out_5_r_bits_id(bus_auto_out_5_r_bits_id),
    .auto_out_5_r_bits_data(bus_auto_out_5_r_bits_data),
    .auto_out_5_r_bits_resp(bus_auto_out_5_r_bits_resp),
    .auto_out_5_r_bits_last(bus_auto_out_5_r_bits_last),
    .auto_out_4_aw_ready(bus_auto_out_4_aw_ready),
    .auto_out_4_aw_valid(bus_auto_out_4_aw_valid),
    .auto_out_4_aw_bits_id(bus_auto_out_4_aw_bits_id),
    .auto_out_4_aw_bits_addr(bus_auto_out_4_aw_bits_addr),
    .auto_out_4_aw_bits_size(bus_auto_out_4_aw_bits_size),
    .auto_out_4_w_ready(bus_auto_out_4_w_ready),
    .auto_out_4_w_valid(bus_auto_out_4_w_valid),
    .auto_out_4_w_bits_data(bus_auto_out_4_w_bits_data),
    .auto_out_4_w_bits_strb(bus_auto_out_4_w_bits_strb),
    .auto_out_4_b_ready(bus_auto_out_4_b_ready),
    .auto_out_4_b_valid(bus_auto_out_4_b_valid),
    .auto_out_4_b_bits_id(bus_auto_out_4_b_bits_id),
    .auto_out_4_b_bits_resp(bus_auto_out_4_b_bits_resp),
    .auto_out_4_ar_ready(bus_auto_out_4_ar_ready),
    .auto_out_4_ar_valid(bus_auto_out_4_ar_valid),
    .auto_out_4_ar_bits_id(bus_auto_out_4_ar_bits_id),
    .auto_out_4_ar_bits_addr(bus_auto_out_4_ar_bits_addr),
    .auto_out_4_ar_bits_size(bus_auto_out_4_ar_bits_size),
    .auto_out_4_r_ready(bus_auto_out_4_r_ready),
    .auto_out_4_r_valid(bus_auto_out_4_r_valid),
    .auto_out_4_r_bits_id(bus_auto_out_4_r_bits_id),
    .auto_out_4_r_bits_data(bus_auto_out_4_r_bits_data),
    .auto_out_4_r_bits_resp(bus_auto_out_4_r_bits_resp),
    .auto_out_4_r_bits_last(bus_auto_out_4_r_bits_last),
    .auto_out_3_aw_ready(bus_auto_out_3_aw_ready),
    .auto_out_3_aw_valid(bus_auto_out_3_aw_valid),
    .auto_out_3_aw_bits_id(bus_auto_out_3_aw_bits_id),
    .auto_out_3_aw_bits_addr(bus_auto_out_3_aw_bits_addr),
    .auto_out_3_aw_bits_size(bus_auto_out_3_aw_bits_size),
    .auto_out_3_w_ready(bus_auto_out_3_w_ready),
    .auto_out_3_w_valid(bus_auto_out_3_w_valid),
    .auto_out_3_w_bits_data(bus_auto_out_3_w_bits_data),
    .auto_out_3_w_bits_strb(bus_auto_out_3_w_bits_strb),
    .auto_out_3_b_ready(bus_auto_out_3_b_ready),
    .auto_out_3_b_valid(bus_auto_out_3_b_valid),
    .auto_out_3_b_bits_id(bus_auto_out_3_b_bits_id),
    .auto_out_3_b_bits_resp(bus_auto_out_3_b_bits_resp),
    .auto_out_3_ar_ready(bus_auto_out_3_ar_ready),
    .auto_out_3_ar_valid(bus_auto_out_3_ar_valid),
    .auto_out_3_ar_bits_id(bus_auto_out_3_ar_bits_id),
    .auto_out_3_ar_bits_addr(bus_auto_out_3_ar_bits_addr),
    .auto_out_3_ar_bits_size(bus_auto_out_3_ar_bits_size),
    .auto_out_3_r_ready(bus_auto_out_3_r_ready),
    .auto_out_3_r_valid(bus_auto_out_3_r_valid),
    .auto_out_3_r_bits_id(bus_auto_out_3_r_bits_id),
    .auto_out_3_r_bits_data(bus_auto_out_3_r_bits_data),
    .auto_out_3_r_bits_resp(bus_auto_out_3_r_bits_resp),
    .auto_out_3_r_bits_last(bus_auto_out_3_r_bits_last),
    .auto_out_2_aw_ready(bus_auto_out_2_aw_ready),
    .auto_out_2_aw_valid(bus_auto_out_2_aw_valid),
    .auto_out_2_aw_bits_id(bus_auto_out_2_aw_bits_id),
    .auto_out_2_aw_bits_addr(bus_auto_out_2_aw_bits_addr),
    .auto_out_2_aw_bits_size(bus_auto_out_2_aw_bits_size),
    .auto_out_2_w_ready(bus_auto_out_2_w_ready),
    .auto_out_2_w_valid(bus_auto_out_2_w_valid),
    .auto_out_2_w_bits_data(bus_auto_out_2_w_bits_data),
    .auto_out_2_w_bits_strb(bus_auto_out_2_w_bits_strb),
    .auto_out_2_b_ready(bus_auto_out_2_b_ready),
    .auto_out_2_b_valid(bus_auto_out_2_b_valid),
    .auto_out_2_b_bits_id(bus_auto_out_2_b_bits_id),
    .auto_out_2_b_bits_resp(bus_auto_out_2_b_bits_resp),
    .auto_out_2_ar_ready(bus_auto_out_2_ar_ready),
    .auto_out_2_ar_valid(bus_auto_out_2_ar_valid),
    .auto_out_2_ar_bits_id(bus_auto_out_2_ar_bits_id),
    .auto_out_2_ar_bits_addr(bus_auto_out_2_ar_bits_addr),
    .auto_out_2_ar_bits_size(bus_auto_out_2_ar_bits_size),
    .auto_out_2_r_ready(bus_auto_out_2_r_ready),
    .auto_out_2_r_valid(bus_auto_out_2_r_valid),
    .auto_out_2_r_bits_id(bus_auto_out_2_r_bits_id),
    .auto_out_2_r_bits_data(bus_auto_out_2_r_bits_data),
    .auto_out_2_r_bits_resp(bus_auto_out_2_r_bits_resp),
    .auto_out_2_r_bits_last(bus_auto_out_2_r_bits_last),
    .auto_out_1_aw_ready(bus_auto_out_1_aw_ready),
    .auto_out_1_aw_valid(bus_auto_out_1_aw_valid),
    .auto_out_1_aw_bits_id(bus_auto_out_1_aw_bits_id),
    .auto_out_1_aw_bits_addr(bus_auto_out_1_aw_bits_addr),
    .auto_out_1_aw_bits_size(bus_auto_out_1_aw_bits_size),
    .auto_out_1_w_ready(bus_auto_out_1_w_ready),
    .auto_out_1_w_valid(bus_auto_out_1_w_valid),
    .auto_out_1_w_bits_data(bus_auto_out_1_w_bits_data),
    .auto_out_1_w_bits_strb(bus_auto_out_1_w_bits_strb),
    .auto_out_1_b_ready(bus_auto_out_1_b_ready),
    .auto_out_1_b_valid(bus_auto_out_1_b_valid),
    .auto_out_1_b_bits_id(bus_auto_out_1_b_bits_id),
    .auto_out_1_b_bits_resp(bus_auto_out_1_b_bits_resp),
    .auto_out_1_ar_ready(bus_auto_out_1_ar_ready),
    .auto_out_1_ar_valid(bus_auto_out_1_ar_valid),
    .auto_out_1_ar_bits_id(bus_auto_out_1_ar_bits_id),
    .auto_out_1_ar_bits_addr(bus_auto_out_1_ar_bits_addr),
    .auto_out_1_ar_bits_size(bus_auto_out_1_ar_bits_size),
    .auto_out_1_r_ready(bus_auto_out_1_r_ready),
    .auto_out_1_r_valid(bus_auto_out_1_r_valid),
    .auto_out_1_r_bits_id(bus_auto_out_1_r_bits_id),
    .auto_out_1_r_bits_data(bus_auto_out_1_r_bits_data),
    .auto_out_1_r_bits_resp(bus_auto_out_1_r_bits_resp),
    .auto_out_1_r_bits_last(bus_auto_out_1_r_bits_last),
    .auto_out_0_aw_ready(bus_auto_out_0_aw_ready),
    .auto_out_0_aw_valid(bus_auto_out_0_aw_valid),
    .auto_out_0_aw_bits_id(bus_auto_out_0_aw_bits_id),
    .auto_out_0_aw_bits_addr(bus_auto_out_0_aw_bits_addr),
    .auto_out_0_aw_bits_size(bus_auto_out_0_aw_bits_size),
    .auto_out_0_w_ready(bus_auto_out_0_w_ready),
    .auto_out_0_w_valid(bus_auto_out_0_w_valid),
    .auto_out_0_w_bits_data(bus_auto_out_0_w_bits_data),
    .auto_out_0_w_bits_strb(bus_auto_out_0_w_bits_strb),
    .auto_out_0_b_ready(bus_auto_out_0_b_ready),
    .auto_out_0_b_valid(bus_auto_out_0_b_valid),
    .auto_out_0_b_bits_id(bus_auto_out_0_b_bits_id),
    .auto_out_0_b_bits_resp(bus_auto_out_0_b_bits_resp),
    .auto_out_0_ar_ready(bus_auto_out_0_ar_ready),
    .auto_out_0_ar_valid(bus_auto_out_0_ar_valid),
    .auto_out_0_ar_bits_id(bus_auto_out_0_ar_bits_id),
    .auto_out_0_ar_bits_addr(bus_auto_out_0_ar_bits_addr),
    .auto_out_0_ar_bits_size(bus_auto_out_0_ar_bits_size),
    .auto_out_0_r_ready(bus_auto_out_0_r_ready),
    .auto_out_0_r_valid(bus_auto_out_0_r_valid),
    .auto_out_0_r_bits_id(bus_auto_out_0_r_bits_id),
    .auto_out_0_r_bits_data(bus_auto_out_0_r_bits_data),
    .auto_out_0_r_bits_resp(bus_auto_out_0_r_bits_resp),
    .auto_out_0_r_bits_last(bus_auto_out_0_r_bits_last)
  );
  AXI4Buffer axi4buf ( // @[Buffer.scala 58:29]
    .clock(axi4buf_clock),
    .reset(axi4buf_reset),
    .auto_in_aw_ready(axi4buf_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_1 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_1_clock),
    .reset(axi4buf_1_reset),
    .auto_in_aw_ready(axi4buf_1_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_1_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_1_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_1_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_1_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_1_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_1_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_1_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_1_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_1_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_1_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_1_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_1_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_1_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_1_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_1_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_1_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_1_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_1_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_1_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_1_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_1_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_1_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_1_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_1_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_1_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_1_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_1_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_1_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_1_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_1_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_1_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_1_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_1_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_1_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_1_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_1_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_1_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_1_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_1_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_1_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_1_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_1_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_1_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_2 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_2_clock),
    .reset(axi4buf_2_reset),
    .auto_in_aw_ready(axi4buf_2_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_2_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_2_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_2_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_2_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_2_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_2_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_2_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_2_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_2_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_2_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_2_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_2_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_2_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_2_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_2_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_2_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_2_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_2_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_2_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_2_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_2_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_2_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_2_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_2_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_2_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_2_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_2_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_2_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_2_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_2_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_2_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_2_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_2_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_2_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_2_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_2_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_2_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_2_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_2_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_2_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_2_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_2_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_2_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_3 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_3_clock),
    .reset(axi4buf_3_reset),
    .auto_in_aw_ready(axi4buf_3_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_3_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_3_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_3_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_3_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_3_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_3_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_3_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_3_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_3_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_3_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_3_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_3_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_3_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_3_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_3_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_3_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_3_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_3_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_3_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_3_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_3_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_3_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_3_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_3_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_3_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_3_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_3_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_3_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_3_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_3_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_3_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_3_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_3_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_3_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_3_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_3_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_3_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_3_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_3_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_3_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_3_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_3_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_3_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_4 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_4_clock),
    .reset(axi4buf_4_reset),
    .auto_in_aw_ready(axi4buf_4_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_4_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_4_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_4_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_4_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_4_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_4_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_4_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_4_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_4_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_4_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_4_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_4_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_4_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_4_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_4_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_4_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_4_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_4_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_4_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_4_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_4_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_4_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_4_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_4_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_4_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_4_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_4_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_4_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_4_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_4_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_4_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_4_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_4_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_4_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_4_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_4_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_4_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_4_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_4_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_4_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_4_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_4_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_4_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_5 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_5_clock),
    .reset(axi4buf_5_reset),
    .auto_in_aw_ready(axi4buf_5_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_5_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_5_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_5_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_5_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_5_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_5_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_5_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_5_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_5_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_5_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_5_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_5_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_5_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_5_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_5_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_5_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_5_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_5_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_5_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_5_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_5_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_5_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_5_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_5_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_5_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_5_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_5_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_5_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_5_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_5_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_5_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_5_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_5_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_5_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_5_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_5_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_5_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_5_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_5_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_5_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_5_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_5_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_5_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_6 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_6_clock),
    .reset(axi4buf_6_reset),
    .auto_in_aw_ready(axi4buf_6_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_6_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_6_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_6_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_6_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_6_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_6_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_6_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_6_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_6_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_6_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_6_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_6_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_6_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_6_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_6_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_6_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_6_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_6_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_6_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_6_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_6_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_6_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_6_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_6_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_6_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_6_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_6_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_6_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_6_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_6_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_6_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_6_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_6_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_6_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_6_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_6_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_6_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_6_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_6_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_6_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_6_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_6_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_6_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_7 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_7_clock),
    .reset(axi4buf_7_reset),
    .auto_in_aw_ready(axi4buf_7_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_7_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_7_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_7_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_7_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_7_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_7_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_7_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_7_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_7_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_7_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_7_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_7_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_7_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_7_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_7_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_7_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_7_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_7_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_7_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_7_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_7_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_7_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_7_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_7_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_7_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_7_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_7_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_7_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_7_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_7_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_7_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_7_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_7_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_7_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_7_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_7_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_7_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_7_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_7_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_7_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_7_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_7_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_7_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_8 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_8_clock),
    .reset(axi4buf_8_reset),
    .auto_in_aw_ready(axi4buf_8_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_8_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_8_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_8_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_8_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_8_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_8_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_8_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_8_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_8_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_8_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_8_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_8_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_8_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_8_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_8_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_8_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_8_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_8_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_8_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_8_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_8_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_8_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_8_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_8_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_8_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_8_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_8_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_8_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_8_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_8_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_8_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_8_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_8_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_8_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_8_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_8_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_8_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_8_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_8_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_8_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_8_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_8_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_8_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_9 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_9_clock),
    .reset(axi4buf_9_reset),
    .auto_in_aw_ready(axi4buf_9_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_9_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_9_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_9_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_9_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_9_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_9_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_9_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_9_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_9_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_9_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_9_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_9_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_9_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_9_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_9_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_9_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_9_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_9_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_9_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_9_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_9_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_9_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_9_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_9_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_9_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_9_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_9_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_9_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_9_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_9_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_9_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_9_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_9_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_9_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_9_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_9_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_9_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_9_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_9_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_9_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_9_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_9_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_9_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_10 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_10_clock),
    .reset(axi4buf_10_reset),
    .auto_in_aw_ready(axi4buf_10_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_10_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_10_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_10_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_10_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_10_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_10_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_10_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_10_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_10_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_10_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_10_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_10_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_10_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_10_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_10_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_10_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_10_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_10_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_10_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_10_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_10_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_10_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_10_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_10_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_10_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_10_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_10_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_10_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_10_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_10_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_10_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_10_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_10_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_10_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_10_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_10_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_10_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_10_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_10_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_10_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_10_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_10_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_10_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_11 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_11_clock),
    .reset(axi4buf_11_reset),
    .auto_in_aw_ready(axi4buf_11_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_11_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_11_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_11_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_11_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_11_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_11_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_11_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_11_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_11_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_11_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_11_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_11_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_11_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_11_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_11_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_11_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_11_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_11_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_11_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_11_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_11_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_11_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_11_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_11_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_11_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_11_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_11_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_11_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_11_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_11_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_11_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_11_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_11_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_11_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_11_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_11_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_11_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_11_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_11_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_11_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_11_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_11_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_11_auto_out_r_bits_data)
  );
  AXI4Buffer axi4buf_12 ( // @[Buffer.scala 58:29]
    .clock(axi4buf_12_clock),
    .reset(axi4buf_12_reset),
    .auto_in_aw_ready(axi4buf_12_auto_in_aw_ready),
    .auto_in_aw_valid(axi4buf_12_auto_in_aw_valid),
    .auto_in_aw_bits_id(axi4buf_12_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(axi4buf_12_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(axi4buf_12_auto_in_aw_bits_size),
    .auto_in_w_ready(axi4buf_12_auto_in_w_ready),
    .auto_in_w_valid(axi4buf_12_auto_in_w_valid),
    .auto_in_w_bits_data(axi4buf_12_auto_in_w_bits_data),
    .auto_in_w_bits_strb(axi4buf_12_auto_in_w_bits_strb),
    .auto_in_b_ready(axi4buf_12_auto_in_b_ready),
    .auto_in_b_valid(axi4buf_12_auto_in_b_valid),
    .auto_in_b_bits_id(axi4buf_12_auto_in_b_bits_id),
    .auto_in_b_bits_resp(axi4buf_12_auto_in_b_bits_resp),
    .auto_in_ar_ready(axi4buf_12_auto_in_ar_ready),
    .auto_in_ar_valid(axi4buf_12_auto_in_ar_valid),
    .auto_in_ar_bits_id(axi4buf_12_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(axi4buf_12_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(axi4buf_12_auto_in_ar_bits_size),
    .auto_in_r_ready(axi4buf_12_auto_in_r_ready),
    .auto_in_r_valid(axi4buf_12_auto_in_r_valid),
    .auto_in_r_bits_id(axi4buf_12_auto_in_r_bits_id),
    .auto_in_r_bits_data(axi4buf_12_auto_in_r_bits_data),
    .auto_in_r_bits_resp(axi4buf_12_auto_in_r_bits_resp),
    .auto_in_r_bits_last(axi4buf_12_auto_in_r_bits_last),
    .auto_out_aw_ready(axi4buf_12_auto_out_aw_ready),
    .auto_out_aw_valid(axi4buf_12_auto_out_aw_valid),
    .auto_out_aw_bits_id(axi4buf_12_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(axi4buf_12_auto_out_aw_bits_addr),
    .auto_out_w_ready(axi4buf_12_auto_out_w_ready),
    .auto_out_w_valid(axi4buf_12_auto_out_w_valid),
    .auto_out_w_bits_data(axi4buf_12_auto_out_w_bits_data),
    .auto_out_w_bits_strb(axi4buf_12_auto_out_w_bits_strb),
    .auto_out_b_ready(axi4buf_12_auto_out_b_ready),
    .auto_out_b_valid(axi4buf_12_auto_out_b_valid),
    .auto_out_b_bits_id(axi4buf_12_auto_out_b_bits_id),
    .auto_out_ar_ready(axi4buf_12_auto_out_ar_ready),
    .auto_out_ar_valid(axi4buf_12_auto_out_ar_valid),
    .auto_out_ar_bits_id(axi4buf_12_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(axi4buf_12_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(axi4buf_12_auto_out_ar_bits_size),
    .auto_out_r_ready(axi4buf_12_auto_out_r_ready),
    .auto_out_r_valid(axi4buf_12_auto_out_r_valid),
    .auto_out_r_bits_id(axi4buf_12_auto_out_r_bits_id),
    .auto_out_r_bits_data(axi4buf_12_auto_out_r_bits_data)
  );
  AXI4StreamBuffer buffer ( // @[Buffer.scala 29:28]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .auto_in_ready(buffer_auto_in_ready),
    .auto_in_valid(buffer_auto_in_valid),
    .auto_in_bits_data(buffer_auto_in_bits_data),
    .auto_in_bits_last(buffer_auto_in_bits_last),
    .auto_out_ready(buffer_auto_out_ready),
    .auto_out_valid(buffer_auto_out_valid),
    .auto_out_bits_data(buffer_auto_out_bits_data),
    .auto_out_bits_last(buffer_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_1 ( // @[Buffer.scala 29:28]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .auto_in_ready(buffer_1_auto_in_ready),
    .auto_in_valid(buffer_1_auto_in_valid),
    .auto_in_bits_data(buffer_1_auto_in_bits_data),
    .auto_in_bits_last(buffer_1_auto_in_bits_last),
    .auto_out_ready(buffer_1_auto_out_ready),
    .auto_out_valid(buffer_1_auto_out_valid),
    .auto_out_bits_data(buffer_1_auto_out_bits_data),
    .auto_out_bits_last(buffer_1_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_2 ( // @[Buffer.scala 29:28]
    .clock(buffer_2_clock),
    .reset(buffer_2_reset),
    .auto_in_ready(buffer_2_auto_in_ready),
    .auto_in_valid(buffer_2_auto_in_valid),
    .auto_in_bits_data(buffer_2_auto_in_bits_data),
    .auto_in_bits_last(buffer_2_auto_in_bits_last),
    .auto_out_ready(buffer_2_auto_out_ready),
    .auto_out_valid(buffer_2_auto_out_valid),
    .auto_out_bits_data(buffer_2_auto_out_bits_data),
    .auto_out_bits_last(buffer_2_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_3 ( // @[Buffer.scala 29:28]
    .clock(buffer_3_clock),
    .reset(buffer_3_reset),
    .auto_in_ready(buffer_3_auto_in_ready),
    .auto_in_valid(buffer_3_auto_in_valid),
    .auto_in_bits_data(buffer_3_auto_in_bits_data),
    .auto_in_bits_last(buffer_3_auto_in_bits_last),
    .auto_out_ready(buffer_3_auto_out_ready),
    .auto_out_valid(buffer_3_auto_out_valid),
    .auto_out_bits_data(buffer_3_auto_out_bits_data),
    .auto_out_bits_last(buffer_3_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_4 ( // @[Buffer.scala 29:28]
    .clock(buffer_4_clock),
    .reset(buffer_4_reset),
    .auto_in_ready(buffer_4_auto_in_ready),
    .auto_in_valid(buffer_4_auto_in_valid),
    .auto_in_bits_data(buffer_4_auto_in_bits_data),
    .auto_in_bits_last(buffer_4_auto_in_bits_last),
    .auto_out_ready(buffer_4_auto_out_ready),
    .auto_out_valid(buffer_4_auto_out_valid),
    .auto_out_bits_data(buffer_4_auto_out_bits_data),
    .auto_out_bits_last(buffer_4_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_5 ( // @[Buffer.scala 29:28]
    .clock(buffer_5_clock),
    .reset(buffer_5_reset),
    .auto_in_ready(buffer_5_auto_in_ready),
    .auto_in_valid(buffer_5_auto_in_valid),
    .auto_in_bits_data(buffer_5_auto_in_bits_data),
    .auto_in_bits_last(buffer_5_auto_in_bits_last),
    .auto_out_ready(buffer_5_auto_out_ready),
    .auto_out_valid(buffer_5_auto_out_valid),
    .auto_out_bits_data(buffer_5_auto_out_bits_data),
    .auto_out_bits_last(buffer_5_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_6 ( // @[Buffer.scala 29:28]
    .clock(buffer_6_clock),
    .reset(buffer_6_reset),
    .auto_in_ready(buffer_6_auto_in_ready),
    .auto_in_valid(buffer_6_auto_in_valid),
    .auto_in_bits_data(buffer_6_auto_in_bits_data),
    .auto_in_bits_last(buffer_6_auto_in_bits_last),
    .auto_out_ready(buffer_6_auto_out_ready),
    .auto_out_valid(buffer_6_auto_out_valid),
    .auto_out_bits_data(buffer_6_auto_out_bits_data),
    .auto_out_bits_last(buffer_6_auto_out_bits_last)
  );
  AXI4StreamBuffer_7 buffer_7 ( // @[Buffer.scala 29:28]
    .clock(buffer_7_clock),
    .reset(buffer_7_reset),
    .auto_in_ready(buffer_7_auto_in_ready),
    .auto_in_valid(buffer_7_auto_in_valid),
    .auto_in_bits_data(buffer_7_auto_in_bits_data),
    .auto_in_bits_last(buffer_7_auto_in_bits_last),
    .auto_out_ready(buffer_7_auto_out_ready),
    .auto_out_valid(buffer_7_auto_out_valid),
    .auto_out_bits_data(buffer_7_auto_out_bits_data),
    .auto_out_bits_last(buffer_7_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_8 ( // @[Buffer.scala 29:28]
    .clock(buffer_8_clock),
    .reset(buffer_8_reset),
    .auto_in_ready(buffer_8_auto_in_ready),
    .auto_in_valid(buffer_8_auto_in_valid),
    .auto_in_bits_data(buffer_8_auto_in_bits_data),
    .auto_in_bits_last(buffer_8_auto_in_bits_last),
    .auto_out_ready(buffer_8_auto_out_ready),
    .auto_out_valid(buffer_8_auto_out_valid),
    .auto_out_bits_data(buffer_8_auto_out_bits_data),
    .auto_out_bits_last(buffer_8_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_9 ( // @[Buffer.scala 29:28]
    .clock(buffer_9_clock),
    .reset(buffer_9_reset),
    .auto_in_ready(buffer_9_auto_in_ready),
    .auto_in_valid(buffer_9_auto_in_valid),
    .auto_in_bits_data(buffer_9_auto_in_bits_data),
    .auto_in_bits_last(buffer_9_auto_in_bits_last),
    .auto_out_ready(buffer_9_auto_out_ready),
    .auto_out_valid(buffer_9_auto_out_valid),
    .auto_out_bits_data(buffer_9_auto_out_bits_data),
    .auto_out_bits_last(buffer_9_auto_out_bits_last)
  );
  AXI4StreamBuffer_7 buffer_10 ( // @[Buffer.scala 29:28]
    .clock(buffer_10_clock),
    .reset(buffer_10_reset),
    .auto_in_ready(buffer_10_auto_in_ready),
    .auto_in_valid(buffer_10_auto_in_valid),
    .auto_in_bits_data(buffer_10_auto_in_bits_data),
    .auto_in_bits_last(buffer_10_auto_in_bits_last),
    .auto_out_ready(buffer_10_auto_out_ready),
    .auto_out_valid(buffer_10_auto_out_valid),
    .auto_out_bits_data(buffer_10_auto_out_bits_data),
    .auto_out_bits_last(buffer_10_auto_out_bits_last)
  );
  AXI4StreamBuffer_7 buffer_11 ( // @[Buffer.scala 29:28]
    .clock(buffer_11_clock),
    .reset(buffer_11_reset),
    .auto_in_ready(buffer_11_auto_in_ready),
    .auto_in_valid(buffer_11_auto_in_valid),
    .auto_in_bits_data(buffer_11_auto_in_bits_data),
    .auto_in_bits_last(buffer_11_auto_in_bits_last),
    .auto_out_ready(buffer_11_auto_out_ready),
    .auto_out_valid(buffer_11_auto_out_valid),
    .auto_out_bits_data(buffer_11_auto_out_bits_data),
    .auto_out_bits_last(buffer_11_auto_out_bits_last)
  );
  AXI4StreamBuffer_7 buffer_12 ( // @[Buffer.scala 29:28]
    .clock(buffer_12_clock),
    .reset(buffer_12_reset),
    .auto_in_ready(buffer_12_auto_in_ready),
    .auto_in_valid(buffer_12_auto_in_valid),
    .auto_in_bits_data(buffer_12_auto_in_bits_data),
    .auto_in_bits_last(buffer_12_auto_in_bits_last),
    .auto_out_ready(buffer_12_auto_out_ready),
    .auto_out_valid(buffer_12_auto_out_valid),
    .auto_out_bits_data(buffer_12_auto_out_bits_data),
    .auto_out_bits_last(buffer_12_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_13 ( // @[Buffer.scala 29:28]
    .clock(buffer_13_clock),
    .reset(buffer_13_reset),
    .auto_in_ready(buffer_13_auto_in_ready),
    .auto_in_valid(buffer_13_auto_in_valid),
    .auto_in_bits_data(buffer_13_auto_in_bits_data),
    .auto_in_bits_last(buffer_13_auto_in_bits_last),
    .auto_out_ready(buffer_13_auto_out_ready),
    .auto_out_valid(buffer_13_auto_out_valid),
    .auto_out_bits_data(buffer_13_auto_out_bits_data),
    .auto_out_bits_last(buffer_13_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_14 ( // @[Buffer.scala 29:28]
    .clock(buffer_14_clock),
    .reset(buffer_14_reset),
    .auto_in_ready(buffer_14_auto_in_ready),
    .auto_in_valid(buffer_14_auto_in_valid),
    .auto_in_bits_data(buffer_14_auto_in_bits_data),
    .auto_in_bits_last(buffer_14_auto_in_bits_last),
    .auto_out_ready(buffer_14_auto_out_ready),
    .auto_out_valid(buffer_14_auto_out_valid),
    .auto_out_bits_data(buffer_14_auto_out_bits_data),
    .auto_out_bits_last(buffer_14_auto_out_bits_last)
  );
  AXI4StreamBuffer buffer_15 ( // @[Buffer.scala 29:28]
    .clock(buffer_15_clock),
    .reset(buffer_15_reset),
    .auto_in_ready(buffer_15_auto_in_ready),
    .auto_in_valid(buffer_15_auto_in_valid),
    .auto_in_bits_data(buffer_15_auto_in_bits_data),
    .auto_in_bits_last(buffer_15_auto_in_bits_last),
    .auto_out_ready(buffer_15_auto_out_ready),
    .auto_out_valid(buffer_15_auto_out_valid),
    .auto_out_bits_data(buffer_15_auto_out_bits_data),
    .auto_out_bits_last(buffer_15_auto_out_bits_last)
  );
  AXI4StreamBuffer_16 buffer_16 ( // @[Buffer.scala 29:28]
    .clock(buffer_16_clock),
    .reset(buffer_16_reset),
    .auto_in_ready(buffer_16_auto_in_ready),
    .auto_in_valid(buffer_16_auto_in_valid),
    .auto_in_bits_data(buffer_16_auto_in_bits_data),
    .auto_in_bits_last(buffer_16_auto_in_bits_last),
    .auto_out_ready(buffer_16_auto_out_ready),
    .auto_out_valid(buffer_16_auto_out_valid),
    .auto_out_bits_data(buffer_16_auto_out_bits_data),
    .auto_out_bits_last(buffer_16_auto_out_bits_last)
  );
  BundleBridgeToAXI4 converter ( // @[Node.scala 65:31]
    .auto_in_aw_ready(converter_auto_in_aw_ready),
    .auto_in_aw_valid(converter_auto_in_aw_valid),
    .auto_in_aw_bits_id(converter_auto_in_aw_bits_id),
    .auto_in_aw_bits_addr(converter_auto_in_aw_bits_addr),
    .auto_in_aw_bits_size(converter_auto_in_aw_bits_size),
    .auto_in_w_ready(converter_auto_in_w_ready),
    .auto_in_w_valid(converter_auto_in_w_valid),
    .auto_in_w_bits_data(converter_auto_in_w_bits_data),
    .auto_in_w_bits_strb(converter_auto_in_w_bits_strb),
    .auto_in_w_bits_last(converter_auto_in_w_bits_last),
    .auto_in_b_ready(converter_auto_in_b_ready),
    .auto_in_b_valid(converter_auto_in_b_valid),
    .auto_in_b_bits_resp(converter_auto_in_b_bits_resp),
    .auto_in_ar_ready(converter_auto_in_ar_ready),
    .auto_in_ar_valid(converter_auto_in_ar_valid),
    .auto_in_ar_bits_id(converter_auto_in_ar_bits_id),
    .auto_in_ar_bits_addr(converter_auto_in_ar_bits_addr),
    .auto_in_ar_bits_size(converter_auto_in_ar_bits_size),
    .auto_in_r_ready(converter_auto_in_r_ready),
    .auto_in_r_valid(converter_auto_in_r_valid),
    .auto_in_r_bits_data(converter_auto_in_r_bits_data),
    .auto_in_r_bits_resp(converter_auto_in_r_bits_resp),
    .auto_in_r_bits_last(converter_auto_in_r_bits_last),
    .auto_out_aw_ready(converter_auto_out_aw_ready),
    .auto_out_aw_valid(converter_auto_out_aw_valid),
    .auto_out_aw_bits_id(converter_auto_out_aw_bits_id),
    .auto_out_aw_bits_addr(converter_auto_out_aw_bits_addr),
    .auto_out_aw_bits_size(converter_auto_out_aw_bits_size),
    .auto_out_w_ready(converter_auto_out_w_ready),
    .auto_out_w_valid(converter_auto_out_w_valid),
    .auto_out_w_bits_data(converter_auto_out_w_bits_data),
    .auto_out_w_bits_strb(converter_auto_out_w_bits_strb),
    .auto_out_w_bits_last(converter_auto_out_w_bits_last),
    .auto_out_b_ready(converter_auto_out_b_ready),
    .auto_out_b_valid(converter_auto_out_b_valid),
    .auto_out_b_bits_resp(converter_auto_out_b_bits_resp),
    .auto_out_ar_ready(converter_auto_out_ar_ready),
    .auto_out_ar_valid(converter_auto_out_ar_valid),
    .auto_out_ar_bits_id(converter_auto_out_ar_bits_id),
    .auto_out_ar_bits_addr(converter_auto_out_ar_bits_addr),
    .auto_out_ar_bits_size(converter_auto_out_ar_bits_size),
    .auto_out_r_ready(converter_auto_out_r_ready),
    .auto_out_r_valid(converter_auto_out_r_valid),
    .auto_out_r_bits_data(converter_auto_out_r_bits_data),
    .auto_out_r_bits_resp(converter_auto_out_r_bits_resp),
    .auto_out_r_bits_last(converter_auto_out_r_bits_last)
  );
  AXI4StreamToBundleBridge converter_1 ( // @[Nodes.scala 165:31]
    .auto_in_ready(converter_1_auto_in_ready),
    .auto_in_valid(converter_1_auto_in_valid),
    .auto_in_bits_data(converter_1_auto_in_bits_data),
    .auto_in_bits_last(converter_1_auto_in_bits_last),
    .auto_out_ready(converter_1_auto_out_ready),
    .auto_out_valid(converter_1_auto_out_valid),
    .auto_out_bits_data(converter_1_auto_out_bits_data),
    .auto_out_bits_last(converter_1_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_2 ( // @[Nodes.scala 201:31]
    .auto_in_ready(converter_2_auto_in_ready),
    .auto_in_valid(converter_2_auto_in_valid),
    .auto_in_bits_data(converter_2_auto_in_bits_data),
    .auto_in_bits_last(converter_2_auto_in_bits_last),
    .auto_out_ready(converter_2_auto_out_ready),
    .auto_out_valid(converter_2_auto_out_valid),
    .auto_out_bits_data(converter_2_auto_out_bits_data),
    .auto_out_bits_last(converter_2_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge_1 converter_3 ( // @[Nodes.scala 165:31]
    .auto_in_ready(converter_3_auto_in_ready),
    .auto_in_valid(converter_3_auto_in_valid),
    .auto_in_bits_data(converter_3_auto_in_bits_data),
    .auto_in_bits_last(converter_3_auto_in_bits_last),
    .auto_out_ready(converter_3_auto_out_ready),
    .auto_out_valid(converter_3_auto_out_valid),
    .auto_out_bits_data(converter_3_auto_out_bits_data),
    .auto_out_bits_last(converter_3_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge_1 converter_4 ( // @[Nodes.scala 165:31]
    .auto_in_ready(converter_4_auto_in_ready),
    .auto_in_valid(converter_4_auto_in_valid),
    .auto_in_bits_data(converter_4_auto_in_bits_data),
    .auto_in_bits_last(converter_4_auto_in_bits_last),
    .auto_out_ready(converter_4_auto_out_ready),
    .auto_out_valid(converter_4_auto_out_valid),
    .auto_out_bits_data(converter_4_auto_out_bits_data),
    .auto_out_bits_last(converter_4_auto_out_bits_last)
  );
  assign ioMem_0_aw_ready = converter_auto_in_aw_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_w_ready = converter_auto_in_w_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_b_valid = converter_auto_in_b_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_b_bits_resp = converter_auto_in_b_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_ar_ready = converter_auto_in_ar_ready; // @[Nodes.scala 624:60]
  assign ioMem_0_r_valid = converter_auto_in_r_valid; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_id = 1'h0; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_data = converter_auto_in_r_bits_data; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_resp = converter_auto_in_r_bits_resp; // @[Nodes.scala 624:60]
  assign ioMem_0_r_bits_last = converter_auto_in_r_bits_last; // @[Nodes.scala 624:60]
  assign outStream_0_valid = converter_1_auto_out_valid; // @[Nodes.scala 649:56]
  assign outStream_0_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign outStream_0_bits_last = converter_1_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign inStream_0_ready = converter_2_auto_in_ready; // @[Nodes.scala 624:60]
  assign laInside_0_valid = converter_3_auto_out_valid; // @[Nodes.scala 649:56]
  assign laInside_0_bits_data = converter_3_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign laInside_0_bits_last = converter_3_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign laOutside_0_valid = converter_4_auto_out_valid; // @[Nodes.scala 649:56]
  assign laOutside_0_bits_data = converter_4_auto_out_bits_data; // @[Nodes.scala 649:56]
  assign laOutside_0_bits_last = converter_4_auto_out_bits_last; // @[Nodes.scala 649:56]
  assign int_0 = uart_int_0; // @[LISTestWithLA.scala 165:9]
  assign uTx = uart_io_txd; // @[LISTestWithLA.scala 171:9]
  assign widthAdapter_clock = clock;
  assign widthAdapter_reset = reset;
  assign widthAdapter_auto_in_valid = in_queue_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_data = in_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_in_bits_last = in_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_auto_out_ready = in_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_clock = clock;
  assign in_split_reset = reset;
  assign in_split_auto_mem_in_aw_valid = axi4buf_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_aw_bits_id = axi4buf_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_aw_bits_addr = axi4buf_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_valid = axi4buf_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_bits_data = axi4buf_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_w_bits_strb = axi4buf_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_b_ready = axi4buf_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_valid = axi4buf_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_id = axi4buf_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_addr = axi4buf_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_ar_bits_size = axi4buf_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign in_split_auto_mem_in_r_ready = axi4buf_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign in_split_auto_stream_in_valid = widthAdapter_auto_out_valid; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_in_bits_data = widthAdapter_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_in_bits_last = widthAdapter_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_4_ready = converter_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_3_ready = buffer_14_auto_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_2_ready = lisFixed_mux0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_1_ready = buffer_3_auto_in_ready; // @[LazyModule.scala 167:57]
  assign in_split_auto_stream_out_0_ready = lisFifo_mux0_auto_stream_in_1_ready; // @[LazyModule.scala 167:57]
  assign in_queue_clock = clock;
  assign in_queue_reset = reset;
  assign in_queue_auto_out_out_ready = widthAdapter_auto_in_ready; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_valid = converter_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_bits_data = converter_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign in_queue_auto_in_in_bits_last = converter_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisFifo_clock = clock;
  assign lisFifo_reset = reset;
  assign lisFifo_auto_mem_in_aw_valid = axi4buf_1_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_aw_bits_id = axi4buf_1_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_aw_bits_addr = axi4buf_1_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_w_valid = axi4buf_1_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_w_bits_data = axi4buf_1_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_w_bits_strb = axi4buf_1_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_b_ready = axi4buf_1_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_ar_valid = axi4buf_1_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_ar_bits_id = axi4buf_1_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_ar_bits_addr = axi4buf_1_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_ar_bits_size = axi4buf_1_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_mem_in_r_ready = axi4buf_1_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_stream_in_valid = lisFifo_mux0_auto_stream_out_0_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_stream_in_bits_data = lisFifo_mux0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_stream_in_bits_last = lisFifo_mux0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:31]
  assign lisFifo_auto_stream_out_ready = buffer_10_auto_in_ready; // @[LazyModule.scala 167:57]
  assign lisFifo_mux0_clock = clock;
  assign lisFifo_mux0_reset = reset;
  assign lisFifo_mux0_auto_register_in_aw_valid = axi4buf_2_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_aw_bits_id = axi4buf_2_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_aw_bits_addr = axi4buf_2_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_w_valid = axi4buf_2_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_w_bits_data = axi4buf_2_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_w_bits_strb = axi4buf_2_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_b_ready = axi4buf_2_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_ar_valid = axi4buf_2_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_ar_bits_id = axi4buf_2_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_ar_bits_addr = axi4buf_2_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_ar_bits_size = axi4buf_2_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_register_in_r_ready = axi4buf_2_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_4_valid = 1'h1; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_4_bits_data = 32'h0; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_4_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_3_valid = 1'h1; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_3_bits_data = 32'hffffffff; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_3_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_2_valid = buffer_1_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_2_bits_data = buffer_1_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_2_bits_last = buffer_1_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_1_valid = in_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign lisFifo_mux0_auto_stream_in_1_bits_data = in_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign lisFifo_mux0_auto_stream_in_1_bits_last = in_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign lisFifo_mux0_auto_stream_in_0_valid = buffer_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_0_bits_data = buffer_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_in_0_bits_last = buffer_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisFifo_mux0_auto_stream_out_0_ready = lisFifo_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign lisInput_clock = clock;
  assign lisInput_reset = reset;
  assign lisInput_auto_mem_in_aw_valid = axi4buf_3_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_aw_bits_id = axi4buf_3_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_aw_bits_addr = axi4buf_3_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_w_valid = axi4buf_3_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_w_bits_data = axi4buf_3_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_w_bits_strb = axi4buf_3_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_b_ready = axi4buf_3_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_ar_valid = axi4buf_3_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_ar_bits_id = axi4buf_3_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_ar_bits_addr = axi4buf_3_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_ar_bits_size = axi4buf_3_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign lisInput_auto_mem_in_r_ready = axi4buf_3_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign lisInput_auto_stream_in_valid = buffer_7_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisInput_auto_stream_in_bits_data = buffer_7_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_auto_stream_in_bits_last = buffer_7_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisInput_auto_stream_out_ready = buffer_11_auto_in_ready; // @[LazyModule.scala 167:57]
  assign lisInput_mux0_clock = clock;
  assign lisInput_mux0_reset = reset;
  assign lisInput_mux0_auto_register_in_aw_valid = axi4buf_4_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_aw_bits_id = axi4buf_4_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_aw_bits_addr = axi4buf_4_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_w_valid = axi4buf_4_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_w_bits_data = axi4buf_4_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_w_bits_strb = axi4buf_4_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_b_ready = axi4buf_4_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_ar_valid = axi4buf_4_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_ar_bits_id = axi4buf_4_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_ar_bits_addr = axi4buf_4_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_ar_bits_size = axi4buf_4_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_register_in_r_ready = axi4buf_4_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_4_valid = buffer_6_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_4_bits_data = buffer_6_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_4_bits_last = buffer_6_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_3_valid = buffer_5_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_3_bits_data = buffer_5_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_3_bits_last = buffer_5_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_2_valid = buffer_4_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_2_bits_data = buffer_4_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_2_bits_last = buffer_4_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_1_valid = buffer_3_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_1_bits_data = buffer_3_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_1_bits_last = buffer_3_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_0_valid = buffer_2_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_0_bits_data = buffer_2_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_in_0_bits_last = buffer_2_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisInput_mux0_auto_stream_out_0_ready = buffer_7_auto_in_ready; // @[LazyModule.scala 167:57]
  assign lisFixed_clock = clock;
  assign lisFixed_reset = reset;
  assign lisFixed_auto_mem_in_aw_valid = axi4buf_5_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_aw_bits_id = axi4buf_5_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_aw_bits_addr = axi4buf_5_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_w_valid = axi4buf_5_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_w_bits_data = axi4buf_5_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_w_bits_strb = axi4buf_5_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_b_ready = axi4buf_5_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_ar_valid = axi4buf_5_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_ar_bits_id = axi4buf_5_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_ar_bits_addr = axi4buf_5_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_ar_bits_size = axi4buf_5_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_mem_in_r_ready = axi4buf_5_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_stream_in_valid = lisFixed_mux0_auto_stream_out_0_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_stream_in_bits_data = lisFixed_mux0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_stream_in_bits_last = lisFixed_mux0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:31]
  assign lisFixed_auto_stream_out_ready = buffer_12_auto_in_ready; // @[LazyModule.scala 167:57]
  assign lisFixed_mux0_clock = clock;
  assign lisFixed_mux0_reset = reset;
  assign lisFixed_mux0_auto_register_in_aw_valid = axi4buf_6_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_aw_bits_id = axi4buf_6_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_aw_bits_addr = axi4buf_6_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_w_valid = axi4buf_6_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_w_bits_data = axi4buf_6_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_w_bits_strb = axi4buf_6_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_b_ready = axi4buf_6_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_ar_valid = axi4buf_6_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_ar_bits_id = axi4buf_6_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_ar_bits_addr = axi4buf_6_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_ar_bits_size = axi4buf_6_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_register_in_r_ready = axi4buf_6_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_4_valid = 1'h1; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_4_bits_data = 32'h0; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_4_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_3_valid = 1'h1; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_3_bits_data = 32'hffffffff; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_3_bits_last = 1'h0; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_2_valid = buffer_9_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_2_bits_data = buffer_9_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_2_bits_last = buffer_9_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_1_valid = in_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:57]
  assign lisFixed_mux0_auto_stream_in_1_bits_data = in_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:57]
  assign lisFixed_mux0_auto_stream_in_1_bits_last = in_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:57]
  assign lisFixed_mux0_auto_stream_in_0_valid = buffer_8_auto_out_valid; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_0_bits_data = buffer_8_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_in_0_bits_last = buffer_8_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign lisFixed_mux0_auto_stream_out_0_ready = lisFixed_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign bist_clock = clock;
  assign bist_reset = reset;
  assign bist_auto_mem_in_aw_valid = axi4buf_7_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_aw_bits_id = axi4buf_7_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_aw_bits_addr = axi4buf_7_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_w_valid = axi4buf_7_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_w_bits_data = axi4buf_7_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_w_bits_strb = axi4buf_7_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_b_ready = axi4buf_7_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_ar_valid = axi4buf_7_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_ar_bits_id = axi4buf_7_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_ar_bits_addr = axi4buf_7_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_ar_bits_size = axi4buf_7_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bist_auto_mem_in_r_ready = axi4buf_7_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bist_auto_stream_out_ready = bist_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign bist_split_clock = clock;
  assign bist_split_reset = reset;
  assign bist_split_auto_mem_in_aw_valid = axi4buf_8_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_aw_bits_id = axi4buf_8_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_aw_bits_addr = axi4buf_8_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_w_valid = axi4buf_8_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_w_bits_data = axi4buf_8_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_w_bits_strb = axi4buf_8_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_b_ready = axi4buf_8_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_ar_valid = axi4buf_8_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_ar_bits_id = axi4buf_8_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_ar_bits_addr = axi4buf_8_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_ar_bits_size = axi4buf_8_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bist_split_auto_mem_in_r_ready = axi4buf_8_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bist_split_auto_stream_in_valid = bist_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign bist_split_auto_stream_in_bits_data = bist_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign bist_split_auto_stream_in_bits_last = bist_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign bist_split_auto_stream_out_3_ready = buffer_13_auto_in_ready; // @[LazyModule.scala 167:57]
  assign bist_split_auto_stream_out_2_ready = buffer_8_auto_in_ready; // @[LazyModule.scala 167:57]
  assign bist_split_auto_stream_out_1_ready = buffer_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign bist_split_auto_stream_out_0_ready = buffer_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_mux_clock = clock;
  assign out_mux_reset = reset;
  assign out_mux_auto_register_in_aw_valid = axi4buf_9_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_aw_bits_id = axi4buf_9_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_aw_bits_addr = axi4buf_9_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_valid = axi4buf_9_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_bits_data = axi4buf_9_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_w_bits_strb = axi4buf_9_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_b_ready = axi4buf_9_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_valid = axi4buf_9_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_id = axi4buf_9_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_addr = axi4buf_9_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_ar_bits_size = axi4buf_9_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign out_mux_auto_register_in_r_ready = axi4buf_9_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_valid = buffer_15_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_bits_data = buffer_15_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_5_bits_last = buffer_15_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_valid = buffer_14_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_bits_data = buffer_14_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_4_bits_last = buffer_14_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_valid = buffer_13_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_bits_data = buffer_13_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_3_bits_last = buffer_13_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_valid = buffer_12_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_bits_data = buffer_12_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_2_bits_last = buffer_12_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_valid = buffer_11_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_bits_data = buffer_11_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_1_bits_last = buffer_11_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_0_valid = buffer_10_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_0_bits_data = buffer_10_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_in_0_bits_last = buffer_10_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_mux_auto_stream_out_1_ready = uTx_queue_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign out_mux_auto_stream_out_0_ready = buffer_16_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_split_clock = clock;
  assign out_split_reset = reset;
  assign out_split_auto_mem_in_aw_valid = axi4buf_10_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_aw_bits_id = axi4buf_10_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_aw_bits_addr = axi4buf_10_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_w_valid = axi4buf_10_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_w_bits_data = axi4buf_10_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_w_bits_strb = axi4buf_10_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_b_ready = axi4buf_10_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_valid = axi4buf_10_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_bits_id = axi4buf_10_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_bits_addr = axi4buf_10_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_ar_bits_size = axi4buf_10_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign out_split_auto_mem_in_r_ready = axi4buf_10_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_in_valid = out_queue_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_in_bits_data = out_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_in_bits_last = out_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:31]
  assign out_split_auto_stream_out_1_ready = converter_4_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_split_auto_stream_out_0_ready = widthAdapter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign out_queue_clock = clock;
  assign out_queue_reset = reset;
  assign out_queue_auto_out_out_ready = out_split_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_valid = buffer_16_auto_out_valid; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_bits_data = buffer_16_auto_out_bits_data; // @[LazyModule.scala 167:31]
  assign out_queue_auto_in_in_bits_last = buffer_16_auto_out_bits_last; // @[LazyModule.scala 167:31]
  assign widthAdapter_1_clock = clock;
  assign widthAdapter_1_reset = reset;
  assign widthAdapter_1_auto_in_valid = out_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_in_bits_data = out_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_in_bits_last = out_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_1_auto_out_ready = converter_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uTx_queue_clock = clock;
  assign uTx_queue_reset = reset;
  assign uTx_queue_auto_out_out_ready = widthAdapter_2_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_valid = out_mux_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_bits_data = out_mux_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign uTx_queue_auto_in_in_bits_last = out_mux_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_clock = clock;
  assign widthAdapter_2_reset = reset;
  assign widthAdapter_2_auto_in_valid = uTx_queue_auto_out_out_valid; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_in_bits_data = uTx_queue_auto_out_out_bits_data; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_in_bits_last = uTx_queue_auto_out_out_bits_last; // @[LazyModule.scala 167:57]
  assign widthAdapter_2_auto_out_ready = uart_auto_in_in_ready; // @[LazyModule.scala 167:57]
  assign widthAdapter_3_clock = clock;
  assign widthAdapter_3_reset = reset;
  assign widthAdapter_3_auto_in_valid = uart_auto_out_out_valid; // @[LazyModule.scala 167:31]
  assign widthAdapter_3_auto_in_bits_data = uart_auto_out_out_bits_data; // @[LazyModule.scala 167:31]
  assign widthAdapter_3_auto_out_ready = uRx_split_auto_stream_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_clock = clock;
  assign uRx_split_reset = reset;
  assign uRx_split_auto_mem_in_aw_valid = axi4buf_12_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_aw_bits_id = axi4buf_12_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_aw_bits_addr = axi4buf_12_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_valid = axi4buf_12_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_bits_data = axi4buf_12_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_w_bits_strb = axi4buf_12_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_b_ready = axi4buf_12_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_valid = axi4buf_12_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_id = axi4buf_12_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_addr = axi4buf_12_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_ar_bits_size = axi4buf_12_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_mem_in_r_ready = axi4buf_12_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign uRx_split_auto_stream_in_valid = widthAdapter_3_auto_out_valid; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_in_bits_data = widthAdapter_3_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_in_bits_last = 1'h0; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_3_ready = buffer_15_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_2_ready = buffer_9_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_1_ready = buffer_4_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uRx_split_auto_stream_out_0_ready = buffer_1_auto_in_ready; // @[LazyModule.scala 167:57]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_auto_mem_in_aw_valid = axi4buf_11_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_aw_bits_id = axi4buf_11_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_aw_bits_addr = axi4buf_11_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_valid = axi4buf_11_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_bits_data = axi4buf_11_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_w_bits_strb = axi4buf_11_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_b_ready = axi4buf_11_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_valid = axi4buf_11_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_id = axi4buf_11_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_addr = axi4buf_11_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_ar_bits_size = axi4buf_11_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign uart_auto_mem_in_r_ready = axi4buf_11_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign uart_auto_in_in_valid = widthAdapter_2_auto_out_valid; // @[LazyModule.scala 167:57]
  assign uart_auto_in_in_bits_data = widthAdapter_2_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign uart_auto_out_out_ready = widthAdapter_3_auto_in_ready; // @[LazyModule.scala 167:31]
  assign uart_io_rxd = uRx; // @[LISTestWithLA.scala 172:24]
  assign bus_clock = clock;
  assign bus_reset = reset;
  assign bus_auto_in_aw_valid = converter_auto_out_aw_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_id = converter_auto_out_aw_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_addr = converter_auto_out_aw_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_aw_bits_size = converter_auto_out_aw_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_valid = converter_auto_out_w_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_data = converter_auto_out_w_bits_data; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_strb = converter_auto_out_w_bits_strb; // @[LazyModule.scala 167:31]
  assign bus_auto_in_w_bits_last = converter_auto_out_w_bits_last; // @[LazyModule.scala 167:31]
  assign bus_auto_in_b_ready = converter_auto_out_b_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_valid = converter_auto_out_ar_valid; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_id = converter_auto_out_ar_bits_id; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_addr = converter_auto_out_ar_bits_addr; // @[LazyModule.scala 167:31]
  assign bus_auto_in_ar_bits_size = converter_auto_out_ar_bits_size; // @[LazyModule.scala 167:31]
  assign bus_auto_in_r_ready = converter_auto_out_r_ready; // @[LazyModule.scala 167:31]
  assign bus_auto_out_12_aw_ready = axi4buf_12_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_w_ready = axi4buf_12_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_valid = axi4buf_12_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_bits_id = axi4buf_12_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_b_bits_resp = axi4buf_12_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_ar_ready = axi4buf_12_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_valid = axi4buf_12_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_id = axi4buf_12_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_data = axi4buf_12_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_resp = axi4buf_12_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_12_r_bits_last = axi4buf_12_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_aw_ready = axi4buf_11_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_w_ready = axi4buf_11_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_valid = axi4buf_11_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_bits_id = axi4buf_11_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_b_bits_resp = axi4buf_11_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_ar_ready = axi4buf_11_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_valid = axi4buf_11_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_id = axi4buf_11_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_data = axi4buf_11_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_resp = axi4buf_11_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_11_r_bits_last = axi4buf_11_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_aw_ready = axi4buf_10_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_w_ready = axi4buf_10_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_valid = axi4buf_10_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_bits_id = axi4buf_10_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_b_bits_resp = axi4buf_10_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_ar_ready = axi4buf_10_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_valid = axi4buf_10_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_id = axi4buf_10_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_data = axi4buf_10_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_resp = axi4buf_10_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_10_r_bits_last = axi4buf_10_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_aw_ready = axi4buf_9_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_w_ready = axi4buf_9_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_valid = axi4buf_9_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_bits_id = axi4buf_9_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_b_bits_resp = axi4buf_9_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_ar_ready = axi4buf_9_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_valid = axi4buf_9_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_id = axi4buf_9_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_data = axi4buf_9_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_resp = axi4buf_9_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_9_r_bits_last = axi4buf_9_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_aw_ready = axi4buf_8_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_w_ready = axi4buf_8_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_valid = axi4buf_8_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_bits_id = axi4buf_8_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_b_bits_resp = axi4buf_8_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_ar_ready = axi4buf_8_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_valid = axi4buf_8_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_id = axi4buf_8_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_data = axi4buf_8_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_resp = axi4buf_8_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_8_r_bits_last = axi4buf_8_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_aw_ready = axi4buf_7_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_w_ready = axi4buf_7_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_valid = axi4buf_7_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_bits_id = axi4buf_7_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_b_bits_resp = axi4buf_7_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_ar_ready = axi4buf_7_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_valid = axi4buf_7_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_id = axi4buf_7_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_data = axi4buf_7_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_resp = axi4buf_7_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_7_r_bits_last = axi4buf_7_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_aw_ready = axi4buf_6_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_w_ready = axi4buf_6_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_valid = axi4buf_6_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_bits_id = axi4buf_6_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_b_bits_resp = axi4buf_6_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_ar_ready = axi4buf_6_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_valid = axi4buf_6_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_id = axi4buf_6_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_data = axi4buf_6_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_resp = axi4buf_6_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_6_r_bits_last = axi4buf_6_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_aw_ready = axi4buf_5_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_w_ready = axi4buf_5_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_valid = axi4buf_5_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_bits_id = axi4buf_5_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_b_bits_resp = axi4buf_5_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_ar_ready = axi4buf_5_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_valid = axi4buf_5_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_id = axi4buf_5_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_data = axi4buf_5_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_resp = axi4buf_5_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_5_r_bits_last = axi4buf_5_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_aw_ready = axi4buf_4_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_w_ready = axi4buf_4_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_valid = axi4buf_4_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_bits_id = axi4buf_4_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_b_bits_resp = axi4buf_4_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_ar_ready = axi4buf_4_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_valid = axi4buf_4_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_id = axi4buf_4_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_data = axi4buf_4_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_resp = axi4buf_4_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_4_r_bits_last = axi4buf_4_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_aw_ready = axi4buf_3_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_w_ready = axi4buf_3_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_valid = axi4buf_3_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_bits_id = axi4buf_3_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_b_bits_resp = axi4buf_3_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_ar_ready = axi4buf_3_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_valid = axi4buf_3_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_id = axi4buf_3_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_data = axi4buf_3_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_resp = axi4buf_3_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_3_r_bits_last = axi4buf_3_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_aw_ready = axi4buf_2_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_w_ready = axi4buf_2_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_valid = axi4buf_2_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_bits_id = axi4buf_2_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_b_bits_resp = axi4buf_2_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_ar_ready = axi4buf_2_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_valid = axi4buf_2_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_id = axi4buf_2_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_data = axi4buf_2_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_resp = axi4buf_2_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_2_r_bits_last = axi4buf_2_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_aw_ready = axi4buf_1_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_w_ready = axi4buf_1_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_valid = axi4buf_1_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_id = axi4buf_1_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_b_bits_resp = axi4buf_1_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_ar_ready = axi4buf_1_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_valid = axi4buf_1_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_id = axi4buf_1_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_data = axi4buf_1_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_resp = axi4buf_1_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_1_r_bits_last = axi4buf_1_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_aw_ready = axi4buf_auto_in_aw_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_w_ready = axi4buf_auto_in_w_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_valid = axi4buf_auto_in_b_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_id = axi4buf_auto_in_b_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_b_bits_resp = axi4buf_auto_in_b_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_ar_ready = axi4buf_auto_in_ar_ready; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_valid = axi4buf_auto_in_r_valid; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_id = axi4buf_auto_in_r_bits_id; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_data = axi4buf_auto_in_r_bits_data; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_resp = axi4buf_auto_in_r_bits_resp; // @[LazyModule.scala 167:57]
  assign bus_auto_out_0_r_bits_last = axi4buf_auto_in_r_bits_last; // @[LazyModule.scala 167:57]
  assign axi4buf_clock = clock;
  assign axi4buf_reset = reset;
  assign axi4buf_auto_in_aw_valid = bus_auto_out_0_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_id = bus_auto_out_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_addr = bus_auto_out_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_aw_bits_size = bus_auto_out_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_valid = bus_auto_out_0_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_data = bus_auto_out_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_w_bits_strb = bus_auto_out_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_b_ready = bus_auto_out_0_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_valid = bus_auto_out_0_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_id = bus_auto_out_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_addr = bus_auto_out_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_ar_bits_size = bus_auto_out_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_in_r_ready = bus_auto_out_0_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_auto_out_aw_ready = in_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_w_ready = in_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_valid = in_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_b_bits_id = in_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_ar_ready = in_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_valid = in_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_id = in_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_auto_out_r_bits_data = in_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_1_clock = clock;
  assign axi4buf_1_reset = reset;
  assign axi4buf_1_auto_in_aw_valid = bus_auto_out_1_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_id = bus_auto_out_1_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_addr = bus_auto_out_1_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_aw_bits_size = bus_auto_out_1_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_valid = bus_auto_out_1_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_data = bus_auto_out_1_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_w_bits_strb = bus_auto_out_1_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_b_ready = bus_auto_out_1_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_valid = bus_auto_out_1_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_id = bus_auto_out_1_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_addr = bus_auto_out_1_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_ar_bits_size = bus_auto_out_1_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_in_r_ready = bus_auto_out_1_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_1_auto_out_aw_ready = lisFifo_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_w_ready = lisFifo_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_valid = lisFifo_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_b_bits_id = lisFifo_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_ar_ready = lisFifo_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_valid = lisFifo_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_id = lisFifo_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_1_auto_out_r_bits_data = lisFifo_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_2_clock = clock;
  assign axi4buf_2_reset = reset;
  assign axi4buf_2_auto_in_aw_valid = bus_auto_out_2_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_id = bus_auto_out_2_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_addr = bus_auto_out_2_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_aw_bits_size = bus_auto_out_2_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_valid = bus_auto_out_2_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_data = bus_auto_out_2_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_w_bits_strb = bus_auto_out_2_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_b_ready = bus_auto_out_2_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_valid = bus_auto_out_2_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_id = bus_auto_out_2_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_addr = bus_auto_out_2_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_ar_bits_size = bus_auto_out_2_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_in_r_ready = bus_auto_out_2_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_2_auto_out_aw_ready = lisFifo_mux0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_w_ready = lisFifo_mux0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_valid = lisFifo_mux0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_b_bits_id = lisFifo_mux0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_ar_ready = lisFifo_mux0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_valid = lisFifo_mux0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_id = lisFifo_mux0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_2_auto_out_r_bits_data = lisFifo_mux0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_3_clock = clock;
  assign axi4buf_3_reset = reset;
  assign axi4buf_3_auto_in_aw_valid = bus_auto_out_3_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_id = bus_auto_out_3_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_addr = bus_auto_out_3_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_aw_bits_size = bus_auto_out_3_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_valid = bus_auto_out_3_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_data = bus_auto_out_3_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_w_bits_strb = bus_auto_out_3_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_b_ready = bus_auto_out_3_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_valid = bus_auto_out_3_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_id = bus_auto_out_3_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_addr = bus_auto_out_3_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_ar_bits_size = bus_auto_out_3_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_in_r_ready = bus_auto_out_3_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_3_auto_out_aw_ready = lisInput_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_w_ready = lisInput_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_valid = lisInput_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_b_bits_id = lisInput_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_ar_ready = lisInput_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_valid = lisInput_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_id = lisInput_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_3_auto_out_r_bits_data = lisInput_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_4_clock = clock;
  assign axi4buf_4_reset = reset;
  assign axi4buf_4_auto_in_aw_valid = bus_auto_out_4_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_id = bus_auto_out_4_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_addr = bus_auto_out_4_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_aw_bits_size = bus_auto_out_4_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_valid = bus_auto_out_4_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_data = bus_auto_out_4_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_w_bits_strb = bus_auto_out_4_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_b_ready = bus_auto_out_4_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_valid = bus_auto_out_4_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_id = bus_auto_out_4_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_addr = bus_auto_out_4_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_ar_bits_size = bus_auto_out_4_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_in_r_ready = bus_auto_out_4_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_4_auto_out_aw_ready = lisInput_mux0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_w_ready = lisInput_mux0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_valid = lisInput_mux0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_b_bits_id = lisInput_mux0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_ar_ready = lisInput_mux0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_valid = lisInput_mux0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_id = lisInput_mux0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_4_auto_out_r_bits_data = lisInput_mux0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_5_clock = clock;
  assign axi4buf_5_reset = reset;
  assign axi4buf_5_auto_in_aw_valid = bus_auto_out_5_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_id = bus_auto_out_5_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_addr = bus_auto_out_5_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_aw_bits_size = bus_auto_out_5_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_valid = bus_auto_out_5_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_data = bus_auto_out_5_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_w_bits_strb = bus_auto_out_5_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_b_ready = bus_auto_out_5_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_valid = bus_auto_out_5_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_id = bus_auto_out_5_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_addr = bus_auto_out_5_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_ar_bits_size = bus_auto_out_5_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_in_r_ready = bus_auto_out_5_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_5_auto_out_aw_ready = lisFixed_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_w_ready = lisFixed_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_valid = lisFixed_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_b_bits_id = lisFixed_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_ar_ready = lisFixed_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_valid = lisFixed_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_id = lisFixed_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_5_auto_out_r_bits_data = lisFixed_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_6_clock = clock;
  assign axi4buf_6_reset = reset;
  assign axi4buf_6_auto_in_aw_valid = bus_auto_out_6_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_id = bus_auto_out_6_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_addr = bus_auto_out_6_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_aw_bits_size = bus_auto_out_6_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_valid = bus_auto_out_6_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_data = bus_auto_out_6_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_w_bits_strb = bus_auto_out_6_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_b_ready = bus_auto_out_6_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_valid = bus_auto_out_6_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_id = bus_auto_out_6_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_addr = bus_auto_out_6_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_ar_bits_size = bus_auto_out_6_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_in_r_ready = bus_auto_out_6_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_6_auto_out_aw_ready = lisFixed_mux0_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_w_ready = lisFixed_mux0_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_valid = lisFixed_mux0_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_b_bits_id = lisFixed_mux0_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_ar_ready = lisFixed_mux0_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_valid = lisFixed_mux0_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_id = lisFixed_mux0_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_6_auto_out_r_bits_data = lisFixed_mux0_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_7_clock = clock;
  assign axi4buf_7_reset = reset;
  assign axi4buf_7_auto_in_aw_valid = bus_auto_out_7_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_id = bus_auto_out_7_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_addr = bus_auto_out_7_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_aw_bits_size = bus_auto_out_7_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_valid = bus_auto_out_7_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_data = bus_auto_out_7_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_w_bits_strb = bus_auto_out_7_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_b_ready = bus_auto_out_7_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_valid = bus_auto_out_7_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_id = bus_auto_out_7_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_addr = bus_auto_out_7_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_ar_bits_size = bus_auto_out_7_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_in_r_ready = bus_auto_out_7_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_7_auto_out_aw_ready = bist_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_w_ready = bist_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_valid = bist_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_b_bits_id = bist_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_ar_ready = bist_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_valid = bist_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_id = bist_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_7_auto_out_r_bits_data = bist_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_8_clock = clock;
  assign axi4buf_8_reset = reset;
  assign axi4buf_8_auto_in_aw_valid = bus_auto_out_8_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_id = bus_auto_out_8_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_addr = bus_auto_out_8_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_aw_bits_size = bus_auto_out_8_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_valid = bus_auto_out_8_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_data = bus_auto_out_8_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_w_bits_strb = bus_auto_out_8_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_b_ready = bus_auto_out_8_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_valid = bus_auto_out_8_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_id = bus_auto_out_8_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_addr = bus_auto_out_8_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_ar_bits_size = bus_auto_out_8_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_in_r_ready = bus_auto_out_8_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_8_auto_out_aw_ready = bist_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_w_ready = bist_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_valid = bist_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_b_bits_id = bist_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_ar_ready = bist_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_valid = bist_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_id = bist_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_8_auto_out_r_bits_data = bist_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_9_clock = clock;
  assign axi4buf_9_reset = reset;
  assign axi4buf_9_auto_in_aw_valid = bus_auto_out_9_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_id = bus_auto_out_9_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_addr = bus_auto_out_9_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_aw_bits_size = bus_auto_out_9_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_valid = bus_auto_out_9_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_data = bus_auto_out_9_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_w_bits_strb = bus_auto_out_9_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_b_ready = bus_auto_out_9_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_valid = bus_auto_out_9_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_id = bus_auto_out_9_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_addr = bus_auto_out_9_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_ar_bits_size = bus_auto_out_9_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_in_r_ready = bus_auto_out_9_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_9_auto_out_aw_ready = out_mux_auto_register_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_w_ready = out_mux_auto_register_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_valid = out_mux_auto_register_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_b_bits_id = out_mux_auto_register_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_ar_ready = out_mux_auto_register_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_valid = out_mux_auto_register_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_id = out_mux_auto_register_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_9_auto_out_r_bits_data = out_mux_auto_register_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_10_clock = clock;
  assign axi4buf_10_reset = reset;
  assign axi4buf_10_auto_in_aw_valid = bus_auto_out_10_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_id = bus_auto_out_10_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_addr = bus_auto_out_10_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_aw_bits_size = bus_auto_out_10_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_valid = bus_auto_out_10_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_data = bus_auto_out_10_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_w_bits_strb = bus_auto_out_10_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_b_ready = bus_auto_out_10_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_valid = bus_auto_out_10_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_id = bus_auto_out_10_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_addr = bus_auto_out_10_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_ar_bits_size = bus_auto_out_10_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_in_r_ready = bus_auto_out_10_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_10_auto_out_aw_ready = out_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_w_ready = out_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_valid = out_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_b_bits_id = out_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_ar_ready = out_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_valid = out_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_id = out_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_10_auto_out_r_bits_data = out_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_11_clock = clock;
  assign axi4buf_11_reset = reset;
  assign axi4buf_11_auto_in_aw_valid = bus_auto_out_11_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_id = bus_auto_out_11_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_addr = bus_auto_out_11_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_aw_bits_size = bus_auto_out_11_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_valid = bus_auto_out_11_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_data = bus_auto_out_11_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_w_bits_strb = bus_auto_out_11_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_b_ready = bus_auto_out_11_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_valid = bus_auto_out_11_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_id = bus_auto_out_11_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_addr = bus_auto_out_11_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_ar_bits_size = bus_auto_out_11_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_in_r_ready = bus_auto_out_11_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_11_auto_out_aw_ready = uart_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_w_ready = uart_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_valid = uart_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_b_bits_id = uart_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_ar_ready = uart_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_valid = uart_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_id = uart_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_11_auto_out_r_bits_data = uart_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign axi4buf_12_clock = clock;
  assign axi4buf_12_reset = reset;
  assign axi4buf_12_auto_in_aw_valid = bus_auto_out_12_aw_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_id = bus_auto_out_12_aw_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_addr = bus_auto_out_12_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_aw_bits_size = bus_auto_out_12_aw_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_valid = bus_auto_out_12_w_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_data = bus_auto_out_12_w_bits_data; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_w_bits_strb = bus_auto_out_12_w_bits_strb; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_b_ready = bus_auto_out_12_b_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_valid = bus_auto_out_12_ar_valid; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_id = bus_auto_out_12_ar_bits_id; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_addr = bus_auto_out_12_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_ar_bits_size = bus_auto_out_12_ar_bits_size; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_in_r_ready = bus_auto_out_12_r_ready; // @[LazyModule.scala 167:57]
  assign axi4buf_12_auto_out_aw_ready = uRx_split_auto_mem_in_aw_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_w_ready = uRx_split_auto_mem_in_w_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_valid = uRx_split_auto_mem_in_b_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_b_bits_id = uRx_split_auto_mem_in_b_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_ar_ready = uRx_split_auto_mem_in_ar_ready; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_valid = uRx_split_auto_mem_in_r_valid; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_id = uRx_split_auto_mem_in_r_bits_id; // @[LazyModule.scala 167:31]
  assign axi4buf_12_auto_out_r_bits_data = uRx_split_auto_mem_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_auto_in_valid = bist_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_data = bist_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_auto_in_bits_last = bist_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_auto_out_ready = lisFifo_mux0_auto_stream_in_0_ready; // @[LazyModule.scala 167:31]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign buffer_1_auto_in_valid = uRx_split_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_data = uRx_split_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_in_bits_last = uRx_split_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_1_auto_out_ready = lisFifo_mux0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign buffer_2_clock = clock;
  assign buffer_2_reset = reset;
  assign buffer_2_auto_in_valid = bist_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_data = bist_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_in_bits_last = bist_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_2_auto_out_ready = lisInput_mux0_auto_stream_in_0_ready; // @[LazyModule.scala 167:31]
  assign buffer_3_clock = clock;
  assign buffer_3_reset = reset;
  assign buffer_3_auto_in_valid = in_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_data = in_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_in_bits_last = in_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_3_auto_out_ready = lisInput_mux0_auto_stream_in_1_ready; // @[LazyModule.scala 167:31]
  assign buffer_4_clock = clock;
  assign buffer_4_reset = reset;
  assign buffer_4_auto_in_valid = uRx_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_in_bits_data = uRx_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_in_bits_last = uRx_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_4_auto_out_ready = lisInput_mux0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign buffer_5_clock = clock;
  assign buffer_5_reset = reset;
  assign buffer_5_auto_in_valid = 1'h1; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_in_bits_data = 32'hffffffff; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_in_bits_last = 1'h0; // @[LazyModule.scala 167:57]
  assign buffer_5_auto_out_ready = lisInput_mux0_auto_stream_in_3_ready; // @[LazyModule.scala 167:31]
  assign buffer_6_clock = clock;
  assign buffer_6_reset = reset;
  assign buffer_6_auto_in_valid = 1'h1; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_in_bits_data = 32'h0; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_in_bits_last = 1'h0; // @[LazyModule.scala 167:57]
  assign buffer_6_auto_out_ready = lisInput_mux0_auto_stream_in_4_ready; // @[LazyModule.scala 167:31]
  assign buffer_7_clock = clock;
  assign buffer_7_reset = reset;
  assign buffer_7_auto_in_valid = lisInput_mux0_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_in_bits_data = lisInput_mux0_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_in_bits_last = lisInput_mux0_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_7_auto_out_ready = lisInput_auto_stream_in_ready; // @[LazyModule.scala 167:31]
  assign buffer_8_clock = clock;
  assign buffer_8_reset = reset;
  assign buffer_8_auto_in_valid = bist_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_in_bits_data = bist_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_in_bits_last = bist_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_8_auto_out_ready = lisFixed_mux0_auto_stream_in_0_ready; // @[LazyModule.scala 167:31]
  assign buffer_9_clock = clock;
  assign buffer_9_reset = reset;
  assign buffer_9_auto_in_valid = uRx_split_auto_stream_out_2_valid; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_in_bits_data = uRx_split_auto_stream_out_2_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_in_bits_last = uRx_split_auto_stream_out_2_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_9_auto_out_ready = lisFixed_mux0_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign buffer_10_clock = clock;
  assign buffer_10_reset = reset;
  assign buffer_10_auto_in_valid = lisFifo_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_10_auto_in_bits_data = lisFifo_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_10_auto_in_bits_last = lisFifo_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_10_auto_out_ready = out_mux_auto_stream_in_0_ready; // @[LazyModule.scala 167:31]
  assign buffer_11_clock = clock;
  assign buffer_11_reset = reset;
  assign buffer_11_auto_in_valid = lisInput_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_11_auto_in_bits_data = lisInput_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_11_auto_in_bits_last = lisInput_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_11_auto_out_ready = out_mux_auto_stream_in_1_ready; // @[LazyModule.scala 167:31]
  assign buffer_12_clock = clock;
  assign buffer_12_reset = reset;
  assign buffer_12_auto_in_valid = lisFixed_auto_stream_out_valid; // @[LazyModule.scala 167:57]
  assign buffer_12_auto_in_bits_data = lisFixed_auto_stream_out_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_12_auto_in_bits_last = lisFixed_auto_stream_out_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_12_auto_out_ready = out_mux_auto_stream_in_2_ready; // @[LazyModule.scala 167:31]
  assign buffer_13_clock = clock;
  assign buffer_13_reset = reset;
  assign buffer_13_auto_in_valid = bist_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:57]
  assign buffer_13_auto_in_bits_data = bist_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_13_auto_in_bits_last = bist_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_13_auto_out_ready = out_mux_auto_stream_in_3_ready; // @[LazyModule.scala 167:31]
  assign buffer_14_clock = clock;
  assign buffer_14_reset = reset;
  assign buffer_14_auto_in_valid = in_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:57]
  assign buffer_14_auto_in_bits_data = in_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_14_auto_in_bits_last = in_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_14_auto_out_ready = out_mux_auto_stream_in_4_ready; // @[LazyModule.scala 167:31]
  assign buffer_15_clock = clock;
  assign buffer_15_reset = reset;
  assign buffer_15_auto_in_valid = uRx_split_auto_stream_out_3_valid; // @[LazyModule.scala 167:57]
  assign buffer_15_auto_in_bits_data = uRx_split_auto_stream_out_3_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_15_auto_in_bits_last = uRx_split_auto_stream_out_3_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_15_auto_out_ready = out_mux_auto_stream_in_5_ready; // @[LazyModule.scala 167:31]
  assign buffer_16_clock = clock;
  assign buffer_16_reset = reset;
  assign buffer_16_auto_in_valid = out_mux_auto_stream_out_0_valid; // @[LazyModule.scala 167:57]
  assign buffer_16_auto_in_bits_data = out_mux_auto_stream_out_0_bits_data; // @[LazyModule.scala 167:57]
  assign buffer_16_auto_in_bits_last = out_mux_auto_stream_out_0_bits_last; // @[LazyModule.scala 167:57]
  assign buffer_16_auto_out_ready = out_queue_auto_in_in_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_in_aw_valid = ioMem_0_aw_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_id = ioMem_0_aw_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_addr = ioMem_0_aw_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_aw_bits_size = ioMem_0_aw_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_valid = ioMem_0_w_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_data = ioMem_0_w_bits_data; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_strb = ioMem_0_w_bits_strb; // @[LazyModule.scala 167:57]
  assign converter_auto_in_w_bits_last = ioMem_0_w_bits_last; // @[LazyModule.scala 167:57]
  assign converter_auto_in_b_ready = ioMem_0_b_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_valid = ioMem_0_ar_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_id = ioMem_0_ar_bits_id; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_addr = ioMem_0_ar_bits_addr; // @[LazyModule.scala 167:57]
  assign converter_auto_in_ar_bits_size = ioMem_0_ar_bits_size; // @[LazyModule.scala 167:57]
  assign converter_auto_in_r_ready = ioMem_0_r_ready; // @[LazyModule.scala 167:57]
  assign converter_auto_out_aw_ready = bus_auto_in_aw_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_w_ready = bus_auto_in_w_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_valid = bus_auto_in_b_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_b_bits_resp = bus_auto_in_b_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_ar_ready = bus_auto_in_ar_ready; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_valid = bus_auto_in_r_valid; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_data = bus_auto_in_r_bits_data; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_resp = bus_auto_in_r_bits_resp; // @[LazyModule.scala 167:31]
  assign converter_auto_out_r_bits_last = bus_auto_in_r_bits_last; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = widthAdapter_1_auto_out_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = widthAdapter_1_auto_out_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = widthAdapter_1_auto_out_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = outStream_0_ready; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = inStream_0_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = inStream_0_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = inStream_0_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = in_queue_auto_in_in_ready; // @[LazyModule.scala 167:31]
  assign converter_3_auto_in_valid = in_split_auto_stream_out_4_valid; // @[LazyModule.scala 167:57]
  assign converter_3_auto_in_bits_data = in_split_auto_stream_out_4_bits_data; // @[LazyModule.scala 167:57]
  assign converter_3_auto_in_bits_last = in_split_auto_stream_out_4_bits_last; // @[LazyModule.scala 167:57]
  assign converter_3_auto_out_ready = laInside_0_ready; // @[LazyModule.scala 167:31]
  assign converter_4_auto_in_valid = out_split_auto_stream_out_1_valid; // @[LazyModule.scala 167:57]
  assign converter_4_auto_in_bits_data = out_split_auto_stream_out_1_bits_data; // @[LazyModule.scala 167:57]
  assign converter_4_auto_in_bits_last = out_split_auto_stream_out_1_bits_last; // @[LazyModule.scala 167:57]
  assign converter_4_auto_out_ready = laOutside_0_ready; // @[LazyModule.scala 167:31]
endmodule
